From pinard@IRO.UMontreal.CA Tue Nov  6 11:43:10 2001
Received: from mercure.IRO.UMontreal.CA (mercure.IRO.UMontreal.CA [132.204.24.67]) by hera.cwi.nl with ESMTP
	id LAA17460 for <Andries.Brouwer@cwi.nl>; Tue, 6 Nov 2001 11:43:09 +0100 (MET)
Received: from trex.iro.umontreal.ca (trex.iro.umontreal.ca [132.204.26.206])
	by mercure.IRO.UMontreal.CA (8.11.4/8.11.1) with ESMTP id fA6Ah7F13588
	for <Andries.Brouwer@cwi.nl>; Tue, 6 Nov 2001 05:43:07 -0500
Received: (from pinard@localhost)
	by trex.iro.umontreal.ca (8.11.4/8.11.1) id fA6Ah7w21029;
	Tue, 6 Nov 2001 05:43:07 -0500
Date: Tue, 6 Nov 2001 05:43:07 -0500
Message-Id: <200111061043.fA6Ah7w21029@trex.iro.umontreal.ca>
From: Translation Project Robot <translation@IRO.UMontreal.CA>
To: Andries.Brouwer@cwi.nl
Subject: Contents of file `kbd-1.06.sv.po'
MIME-Version: 1.0
Content-Type: multipart/mixed; boundary="=-=-="
Status: R

--=-=-=
Content-Type: application/octet-stream
Content-Disposition: attachment; filename=kbd-1.06.sv.po
Content-Transfer-Encoding: base64

IyBTd2VkaXNoIG1lc3NhZ2UgZmlsZSBmb3Iga2JkCiMgQ29weXJpZ2h0IChDKSAyMDAxIEZyZWUg
U29mdHdhcmUgRm91bmRhdGlvbiwgSW5jLgojIE1hcnRpbiBTavZncmVuIDxtZDltc0BtZHN0dWQu
Y2hhbG1lcnMuc2U+LCAyMDAxLgojCiMgJElkOiBzdi5wbyx2IDEuMTUgMjAwMS8xMS8wNiAxMDoz
NDozMyBtYXJ0aW4gRXhwICQKIwptc2dpZCAiIgptc2dzdHIgIiIKIlByb2plY3QtSWQtVmVyc2lv
bjoga2JkIDEuMDZcbiIKIlBPVC1DcmVhdGlvbi1EYXRlOiAyMDAxLTA5LTMwIDExOjI5KzAyMDBc
biIKIlBPLVJldmlzaW9uLURhdGU6IDIwMDEtMTEtMDYgMTE6MzMrMDEwMFxuIgoiTGFzdC1UcmFu
c2xhdG9yOiBNYXJ0aW4gU2r2Z3JlbiA8bWQ5bXNAbWRzdHVkLmNoYWxtZXJzLnNlPlxuIgoiTGFu
Z3VhZ2UtVGVhbTogU3dlZGlzaCA8c3ZAbGkub3JnPlxuIgoiTUlNRS1WZXJzaW9uOiAxLjBcbiIK
IkNvbnRlbnQtVHlwZTogdGV4dC9wbGFpbjsgY2hhcnNldD1pc28tODg1OS0xXG4iCiJDb250ZW50
LVRyYW5zZmVyLUVuY29kaW5nOiA4Yml0XG4iCgojOiBvcGVudnQvb3BlbnZ0LmM6NjcKIywgYy1m
b3JtYXQKbXNnaWQgIm9wZW52dDogJXM6IGlsbGVnYWwgdnQgbnVtYmVyXG4iCm1zZ3N0ciAib3Bl
bnZ0OiAlczogb2dpbHRpZ3QgdnQtbnVtbWVyXG4iCgojOiBvcGVudnQvb3BlbnZ0LmM6OTEKbXNn
aWQgIm9wZW52dDogb25seSByb290IGNhbiB1c2UgdGhlIC11IGZsYWcuXG4iCm1zZ3N0ciAib3Bl
bnZ0OiBlbmRhc3Qgcm9vdCBrYW4gYW525G5kYSBmbGFnZ2FuIC11LlxuIgoKIzogb3BlbnZ0L29w
ZW52dC5jOjEwNSBzcmMvZ2V0ZmQuYzo2Mwptc2dpZCAiQ291bGRudCBnZXQgYSBmaWxlIGRlc2Ny
aXB0b3IgcmVmZXJyaW5nIHRvIHRoZSBjb25zb2xlXG4iCm1zZ3N0ciAiS3VuZGUgaW50ZSBm5SBl
biBmaWxpZGVudGlmaWVyYXJlIGb2ciBrb25zb2xsZW5cbiIKCiM6IG9wZW52dC9vcGVudnQuYzox
MTcKbXNnaWQgIm9wZW52dDogY2Fubm90IGZpbmQgYSBmcmVlIHZ0XG4iCm1zZ3N0ciAib3BlbnZ0
OiBrYW4gaW50ZSBoaXR0YSBlbiBsZWRpZyB2dFxuIgoKIzogb3BlbnZ0L29wZW52dC5jOjEyMgoj
LCBjLWZvcm1hdAptc2dpZCAib3BlbnZ0OiBjYW5ub3QgY2hlY2sgd2hldGhlciB2dCAlZCBpcyBm
cmVlXG4iCm1zZ3N0ciAib3BlbnZ0OiBrYW4gaW50ZSB1bmRlcnP2a2EgaHVydXZpZGEgdnQgJWQg
5HIgbGVkaWdcbiIKCiM6IG9wZW52dC9vcGVudnQuYzoxMjMgb3BlbnZ0L29wZW52dC5jOjEyOApt
c2dpZCAiICAgICAgICB1c2UgYG9wZW52dCAtZicgdG8gZm9yY2UuXG4iCm1zZ3N0ciAiICAgICAg
ICBhbnbkbmQgXCJvcGVudnQgLWZcIiBm9nIgYXR0IHR2aW5nYS5cbiIKCiM6IG9wZW52dC9vcGVu
dnQuYzoxMjcKIywgYy1mb3JtYXQKbXNnaWQgIm9wZW52dDogdnQgJWQgaXMgaW4gdXNlOyBjb21t
YW5kIGFib3J0ZWRcbiIKbXNnc3RyICJvcGVudnQ6IHZ0ICVkIGFuduRuZHMsIGtvbW1hbmRvdCBh
dmJydXRldFxuIgoKIzogb3BlbnZ0L29wZW52dC5jOjE1NQojLCBjLWZvcm1hdAptc2dpZCAib3Bl
bnZ0OiBVbmFibGUgdG8gb3BlbiAlczogJXNcbiIKbXNnc3RyICJvcGVudnQ6IEthbiBpbnRlIPZw
cG5hICVzOiAlc1xuIgoKIzogb3BlbnZ0L29wZW52dC5jOjE2NwojLCBjLWZvcm1hdAptc2dpZCAi
b3BlbnZ0OiBDYW5ub3Qgb3BlbiAlcyByZWFkL3dyaXRlICglcylcbiIKbXNnc3RyICJvcGVudnQ6
IEthbiBpbnRlIPZwcG5hICVzIGb2ciBs5HNuaW5nL3Nrcml2bmluZyAoJXMpXG4iCgojOiBvcGVu
dnQvb3BlbnZ0LmM6MjA1CiMsIGMtZm9ybWF0Cm1zZ2lkICJvcGVudnQ6IHVzaW5nIFZUICVzXG4i
Cm1zZ3N0ciAib3BlbnZ0OiBhbnbkbmRlciBWVCAlc1xuIgoKIzogb3BlbnZ0L29wZW52dC5jOjIx
NwojLCBjLWZvcm1hdAptc2dpZCAib3BlbnZ0OiBVbmFibGUgdG8gc2V0IG5ldyBzZXNzaW9uICgl
cylcbiIKbXNnc3RyICJvcGVudnQ6IEthbiBpbnRlIHPkdHRhIG55IHNlc3Npb24gKCVzKVxuIgoK
Izogb3BlbnZ0L29wZW52dC5jOjIyNQojLCBjLWZvcm1hdAptc2dpZCAiXG5vcGVudnQ6IGNvdWxk
IG5vdCBvcGVuICVzIFIvVyAoJXMpXG4iCm1zZ3N0ciAiXG5vcGVudnQ6IGt1bmRlIGludGUg9nBw
bmEgJXMgZvZyIGzkc25pbmcvc2tyaXZuaW5nICglcylcbiIKCiM6IG9wZW52dC9vcGVudnQuYzoy
ODEKIywgYy1mb3JtYXQKbXNnaWQgIm9wZW52dDogY291bGQgbm90IGRlYWxsb2NhdGUgY29uc29s
ZSAlZFxuIgptc2dzdHIgIm9wZW52dDoga3VuZGUgaW50ZSBkZWFsbG9rZXJhIGtvbnNvbGwgJWRc
biIKCiM6IHNyYy9jaHZ0LmM6MjgKbXNnaWQgInVzYWdlOiBjaHZ0IE5cbiIKbXNnc3RyICJhbnbk
bmRuaW5nOiBjaHZ0IE5cbiIKCiM6IHNyYy9kZWFsbG9jdnQuYzozMwojLCBjLWZvcm1hdAptc2dp
ZCAiJXM6IHVua25vd24gb3B0aW9uXG4iCm1zZ3N0ciAiJXM6IG9r5G5kIGZsYWdnYVxuIgoKIzog
c3JjL2RlYWxsb2N2dC5jOjQ1CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogZGVhbGxvY2F0aW5nIGFs
bCB1bnVzZWQgY29uc29sZXMgZmFpbGVkXG4iCm1zZ3N0ciAiJXM6IGRlYWxsb2tlcmluZyBhdiBh
bGxhIG9hbnbkbmRhIGtvbnNvbGxlciBtaXNzbHlja2FkZXNcbiIKCiM6IHNyYy9kZWFsbG9jdnQu
Yzo1MwojLCBjLWZvcm1hdAptc2dpZCAiJXM6IDA6IGlsbGVnYWwgVlQgbnVtYmVyXG4iCm1zZ3N0
ciAiJXM6IDA6IG9naWx0aWd0IFZULW51bW1lclxuIgoKIzogc3JjL2RlYWxsb2N2dC5jOjU2CiMs
IGMtZm9ybWF0Cm1zZ2lkICIlczogVlQgMSBpcyB0aGUgY29uc29sZSBhbmQgY2Fubm90IGJlIGRl
YWxsb2NhdGVkXG4iCm1zZ3N0ciAiJXM6IFZUIDEg5HIga29uc29sbGVuIG9jaCBrYW4gaW50ZSBk
ZWFsbG9rZXJhc1xuIgoKIzogc3JjL2RlYWxsb2N2dC5jOjYxCiMsIGMtZm9ybWF0Cm1zZ2lkICIl
czogY291bGQgbm90IGRlYWxsb2NhdGUgY29uc29sZSAlZFxuIgptc2dzdHIgIiVzOiBrdW5kZSBp
bnRlIGRlYWxsb2tlcmEga29uc29sbCAlZFxuIgoKIzogc3JjL2R1bXBrZXlzLmM6NjMKIywgYy1m
b3JtYXQKbXNnaWQgIktER0tCRU5UIGVycm9yIGF0IGluZGV4IDAgaW4gdGFibGUgJWQ6ICIKbXNn
c3RyICJLREdLQkVOVC1mZWwgdmlkIGluZGV4IDAgaSB0YWJlbGwgJWQ6ICIKCiM6IHNyYy9kdW1w
a2V5cy5jOjc2CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogY2Fubm90IGZpbmQgYW55IGtleW1hcHM/
XG4iCm1zZ3N0ciAiJXM6IGthbiBpbnRlIGhpdHRhIG7lZ3JhIHRhbmdlbnR0YWJlbGxlcj9cbiIK
CiM6IHNyYy9kdW1wa2V5cy5jOjgxCiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogcGxhaW4gbWFwIG5v
dCBhbGxvY2F0ZWQ/IHZlcnkgc3RyYW5nZSAuLi5cbiIKbXNnc3RyICIlczogZW5rZWwgdGFiZWxs
IGludGUgYWxsb2tlcmFkPyBteWNrZXQgbXlzdGlza3QgLi4uXG4iCgojOiBzcmMvZHVtcGtleXMu
YzoxMTMKIywgYy1mb3JtYXQKbXNnaWQgIktER0tCRU5UIGVycm9yIGF0IGluZGV4ICVkIGluIHRh
YmxlICVkOiAiCm1zZ3N0ciAiS0RHS0JFTlQtZmVsIHZpZCBpbmRleCAlZCBpIHRhYmVsbCAlZDog
IgoKIzogc3JjL2R1bXBrZXlzLmM6MjQxCiMsIGMtZm9ybWF0Cm1zZ2lkICJrZXljb2RlIHJhbmdl
IHN1cHBvcnRlZCBieSBrZXJuZWw6ICAgICAgICAgICAxIC0gJWRcbiIKbXNnc3RyICJ0YW5nZW50
a29kc2ludGVydmFsbCBzb20gc3T2ZHMgYXYga+RybmFuOiAgICAgICAgMSAtICVkXG4iCgojOiBz
cmMvZHVtcGtleXMuYzoyNDMKIywgYy1mb3JtYXQKbXNnaWQgIm1heCBudW1iZXIgb2YgYWN0aW9u
cyBiaW5kYWJsZSB0byBhIGtleTogICAgICAgICAlZFxuIgptc2dzdHIgInN09nJzdGEgYW50YWwg
aGFuZGxpbmdhciBiaW5kYmFyYSB0aWxsIGVuIHRhbmdlbnQ6ICAgJWRcbiIKCiM6IHNyYy9kdW1w
a2V5cy5jOjI0NgojLCBjLWZvcm1hdAptc2dpZCAibnVtYmVyIG9mIGtleW1hcHMgaW4gYWN0dWFs
IHVzZTogICAgICAgICAgICAgICAgICVkXG4iCm1zZ3N0ciAiYW50YWwgdGFuZ2VudHRhYmVsbGVy
IHNvbSBmYWt0aXNrdCBhbnbkbmRzOiAgICAgICAgICAlZFxuIgoKIzogc3JjL2R1bXBrZXlzLmM6
MjQ5CiMsIGMtZm9ybWF0Cm1zZ2lkICJvZiB3aGljaCAlZCBkeW5hbWljYWxseSBhbGxvY2F0ZWRc
biIKbXNnc3RyICJ2YXJhdiAlZCDkciBkeW5hbWlza3QgYWxsb2tlcmFkZVxuIgoKIzogc3JjL2R1
bXBrZXlzLmM6MjUwCm1zZ2lkICJyYW5nZXMgb2YgYWN0aW9uIGNvZGVzIHN1cHBvcnRlZCBieSBr
ZXJuZWw6XG4iCm1zZ3N0ciAiaW50ZXJ2YWxsIGF2IGhhbmRsaW5nc2tvZGVyIHNvbSBzdPZkcyBh
diBr5HJuYW46XG4iCgojOiBzcmMvZHVtcGtleXMuYzoyNTUKIywgYy1mb3JtYXQKbXNnaWQgIm51
bWJlciBvZiBmdW5jdGlvbiBrZXlzIHN1cHBvcnRlZCBieSBrZXJuZWw6ICVkXG4iCm1zZ3N0ciAi
YW50YWwgZnVua3Rpb25zdGFuZ2VudGVyIHNvbSBzdPZkcyBhdiBr5HJuYW46ICVkXG4iCgojOiBz
cmMvZHVtcGtleXMuYzoyNTgKIywgYy1mb3JtYXQKbXNnaWQgIm1heCBuciBvZiBjb21wb3NlIGRl
ZmluaXRpb25zOiAlZFxuIgptc2dzdHIgInN09nJzdGEgYW50YWwga29tcG9zaXRpb25zZGVmaW5p
dGlvbmVyOiAlZFxuIgoKIzogc3JjL2R1bXBrZXlzLmM6MjYwCiMsIGMtZm9ybWF0Cm1zZ2lkICJu
ciBvZiBjb21wb3NlIGRlZmluaXRpb25zIGluIGFjdHVhbCB1c2U6ICVkXG4iCm1zZ3N0ciAiYW50
YWwga29tcG9zaXRpb25zZGVmaW5pdGlvbmVyIHNvbSBmYWt0aXNrdCBhbnbkbmRzOiAlZFxuIgoK
Izogc3JjL2R1bXBrZXlzLmM6Mjg0CiMsIGMtZm9ybWF0Cm1zZ2lkICIiCiJTeW1ib2xzIHJlY29n
bml6ZWQgYnkgJXM6XG4iCiIobnVtZXJpYyB2YWx1ZSwgc3ltYm9sKVxuIgoiXG4iCm1zZ3N0ciAi
IgoiU3ltYm9sZXIgc29tIGvkbm5zIGlnZW4gYXYgJXM6XG4iCiIobnVtZXJpc2t0IHbkcmRlLCBz
eW1ib2wpXG4iCiJcbiIKCiM6IHNyYy9kdW1wa2V5cy5jOjI5Nwptc2dpZCAiXG5UaGUgZm9sbG93
aW5nIHN5bm9ueW1zIGFyZSByZWNvZ25pemVkOlxuXG4iCm1zZ3N0ciAiXG5G9mxqYW5kZSBzeW5v
bnltZXIga+RubnMgaWdlbjpcblxuIgoKIzogc3JjL2R1bXBrZXlzLmM6Mjk5CiMsIGMtZm9ybWF0
Cm1zZ2lkICIlLTE1cyBmb3IgJXNcbiIKbXNnc3RyICIlLTE1cyBm9nIgJXNcbiIKCiM6IHNyYy9k
dW1wa2V5cy5jOjMwMQptc2dpZCAiXG5SZWNvZ25pemVkIG1vZGlmaWVyIG5hbWVzIGFuZCB0aGVp
ciBjb2x1bW4gbnVtYmVyczpcbiIKbXNnc3RyICJcbklnZW5r5G5kYSBtb2RpZmllcmFybmFtbiBv
Y2ggZGVyYXMga29sdW1ubnVtbWVyOlxuIgoKIzogc3JjL2R1bXBrZXlzLmM6MzY0CiMsIGMtZm9y
bWF0Cm1zZ2lkICIjIG5vdCBhbHRfaXNfbWV0YTogb24ga2V5bWFwICVkIGtleSAlZCBpcyBib3Vu
ZCB0byIKbXNnc3RyICIjIGludGUgYWx0X2lzX21ldGE6IGkgdGFuZ2VudHRhYmVsbCAlZCDkciB0
YW5nZW50ICVkIGJ1bmRlbiB0aWxsIgoKIzogc3JjL2R1bXBrZXlzLmM6NDM5Cm1zZ2lkICJpbXBv
c3NpYmxlOiBub3QgbWV0YT9cbiIKbXNnc3RyICJvbfZqbGlndDogaW50ZSBtZXRhP1xuIgoKIzog
c3JjL2R1bXBrZXlzLmM6NDk2CiMsIGMtZm9ybWF0Cm1zZ2lkICJLREdLQlNFTlQgZmFpbGVkIGF0
IGluZGV4ICVkOiAiCm1zZ3N0ciAiS0RHS0JTRU5UIG1pc3NseWNrYWRlcyB2aWQgaW5kZXggJWQ6
ICIKCiM6IHNyYy9kdW1wa2V5cy5jOjUxNgojLCBjLWZvcm1hdAptc2dpZCAiZHVtcGtleXMgdmVy
c2lvbiAlcyIKbXNnc3RyICJkdW1wa2V5cyB2ZXJzaW9uICVzIgoKIzogc3JjL2R1bXBrZXlzLmM6
NTE3Cm1zZ2lkICIiCiJcbiIKInVzYWdlOiBkdW1wa2V5cyBbb3B0aW9ucy4uLl1cbiIKIlxuIgoi
dmFsaWQgb3B0aW9ucyBhcmU6XG4iCiJcbiIKIlx0LWggLS1oZWxwXHQgICAgZGlzcGxheSB0aGlz
IGhlbHAgdGV4dFxuIgoiXHQtaSAtLXNob3J0LWluZm9cdCAgICBkaXNwbGF5IGluZm9ybWF0aW9u
IGFib3V0IGtleWJvYXJkIGRyaXZlclxuIgoiXHQtbCAtLWxvbmctaW5mb1x0ICAgIGRpc3BsYXkg
YWJvdmUgYW5kIHN5bWJvbHMga25vd24gdG8gbG9hZGtleXNcbiIKIlx0LW4gLS1udW1lcmljXHQg
ICAgZGlzcGxheSBrZXl0YWJsZSBpbiBoZXhhZGVjaW1hbCBub3RhdGlvblxuIgoiXHQtZiAtLWZ1
bGwtdGFibGVcdCAgICBkb24ndCB1c2Ugc2hvcnQtaGFuZCBub3RhdGlvbnMsIG9uZSByb3cgcGVy
IGtleWNvZGVcbiIKIlx0LTEgLS1zZXBhcmF0ZS1saW5lcyBvbmUgbGluZSBwZXIgKG1vZGlmaWVy
LGtleWNvZGUpIHBhaXJcbiIKIlx0ICAgLS1mdW5jcy1vbmx5XHQgICAgZGlzcGxheSBvbmx5IHRo
ZSBmdW5jdGlvbiBrZXkgc3RyaW5nc1xuIgoiXHQgICAtLWtleXMtb25seVx0ICAgIGRpc3BsYXkg
b25seSBrZXkgYmluZGluZ3NcbiIKIlx0ICAgLS1jb21wb3NlLW9ubHkgICBkaXNwbGF5IG9ubHkg
Y29tcG9zZSBrZXkgY29tYmluYXRpb25zXG4iCiJcdC1jIC0tY2hhcnNldD0iCm1zZ3N0ciAiIgoi
XG4iCiJhbnbkbmRuaW5nOiBkdW1wa2V5cyBbZmxhZ2dvci4uLl1cbiIKIlxuIgoiZ2lsdGlnYSBm
bGFnZ29yIORyOlxuIgoiXG4iCiJcdC1oIC0taGVscFx0ICAgIHZpc2EgZGVuIGjkciBoauRscHRl
eHRlblxuIgoiXHQtaSAtLXNob3J0LWluZm9cdCAgICB2aXNhIGluZm9ybWF0aW9uIG9tIHRhbmdl
bnRib3Jkc2RyaXZ1dGluXG4iCiJcdC1sIC0tbG9uZy1pbmZvXHQgICAgdmlzYSBvdmFuc3TlZW5k
ZSBvY2ggc3ltYm9sZXIga+RuZGEgZvZyIGxvYWRrZXlzXG4iCiJcdC1uIC0tbnVtZXJpY1x0ICAg
IHZpc2EgdGFuZ2VudHRhYmVsbCBpIGhleGFkZWNpbWFsIG5vdGF0aW9uXG4iCiJcdC1mIC0tZnVs
bC10YWJsZVx0ICAgIGFuduRuZCBpbnRlIGtvcnQgbm90YXRpb24sIGVuIHJhZCBwZXIgdGFuZ2Vu
dGtvZFxuIgoiXHQtMSAtLXNlcGFyYXRlLWxpbmVzIGVuIHJhZCBwZXIgKG1vZGlmaWVyYXJlLHRh
bmdlbnRrb2QpLXBhclxuIgoiXHQgICAtLWZ1bmNzLW9ubHlcdCAgICB2aXNhIGJhcmEgc3Ry5G5n
YXIgZvZyIGZ1bmt0aW9uc3RhbmdlbnRlclxuIgoiXHQgICAtLWtleXMtb25seVx0ICAgIHZpc2Eg
YmFyYSB0YW5nZW50YmluZG5pbmdhclxuIgoiXHQgICAtLWNvbXBvc2Wtb25seSAgIHZpc2EgYmFy
YSBcImNvbXBvc2VcIi10YW5nZW50a29tYmluYXRpb25lclxuIgoiXHQtYyAtLWNoYXJzZXQ9IgoK
Izogc3JjL2R1bXBrZXlzLmM6NTM0Cm1zZ2lkICIiCiJcdFx0XHQgICAgaW50ZXJwcmV0IGNoYXJh
Y3RlciBhY3Rpb24gY29kZXMgdG8gYmUgZnJvbSB0aGVcbiIKIlx0XHRcdCAgICBzcGVjaWZpZWQg
Y2hhcmFjdGVyIHNldFxuIgptc2dzdHIgIiIKIlx0XHRcdCAgICB0b2xrYSB0ZWNrZW5oYW5kbGlu
Z3Nrb2RlciBzb20gb20gZGUg5HIgZnLlbiBkZW5cbiIKIlx0XHRcdCAgICBhbmdpdm5hIHRlY2tl
bnVwcHPkdHRuaW5nZW5cbiIKCiM6IHNyYy9maW5kZmlsZS5jOjQzCiMsIGMtZm9ybWF0Cm1zZ2lk
ICJlcnJvciBleGVjdXRpbmcgICVzXG4iCm1zZ3N0ciAiZmVsIHZpZCBleGVrdmVyaW5nIGF2ICVz
XG4iCgojOiBzcmMvZ2V0a2V5Y29kZXMuYzoxOAptc2dpZCAidXNhZ2U6IGdldGtleWNvZGVzXG4i
Cm1zZ3N0ciAiYW525G5kbmluZzogZ2V0a2V5Y29kZXNcbiIKCiM6IHNyYy9nZXRrZXljb2Rlcy5j
OjM5Cm1zZ2lkICJQbGFpbiBzY2FuY29kZXMgeHggKGhleCkgdmVyc3VzIGtleWNvZGVzIChkZWMp
XG4iCm1zZ3N0ciAiRW5rbGEgYXZs5HNuaW5nc2tvZGVyIHh4IChoZXgpIG1vdCB0YW5nZW50a29k
ZXIgKGRlYylcbiIKCiM6IHNyYy9nZXRrZXljb2Rlcy5jOjQwCm1zZ2lkICIwIGlzIGFuIGVycm9y
OyBmb3IgMS04OCAoMHgwMS0weDU4KSBzY2FuY29kZSBlcXVhbHMga2V5Y29kZVxuIgptc2dzdHIg
IjAg5HIgZXR0IGZlbCwgZvZyIDEtODggKDB4MDEtMHg1OCkg5HIgYXZs5HNuaW5nc2tvZGVuIGxp
a2EgbWVkIHRhbmdlbnRrb2RlblxuIgoKIzogc3JjL2dldGtleWNvZGVzLmM6NDQKbXNnaWQgIlxu
XG5Fc2NhcGVkIHNjYW5jb2RlcyBlMCB4eCAoaGV4KVxuIgptc2dzdHIgIlxuXG5VdHZpZGdhZGUg
YXZs5HNuaW5nc2tvZGVyIGUwIHh4IChoZXgpXG4iCgojOiBzcmMvZ2V0a2V5Y29kZXMuYzo2NAoj
LCBjLWZvcm1hdAptc2dpZCAiZmFpbGVkIHRvIGdldCBrZXljb2RlIGZvciBzY2FuY29kZSAweCV4
XG4iCm1zZ3N0ciAibWlzc2x5Y2thZGVzIG1lZCBhdHQgaORtdGEgdGFuZ2VudGtvZGVuIGb2ciBh
dmzkc25pbmdza29kIDB4JXhcbiIKCiM6IHNyYy9nZXR1bmltYXAuYzo0OQojLCBjLWZvcm1hdApt
c2dpZCAiIgoiVXNhZ2U6XG4iCiJcdCVzIFstc11cbiIKbXNnc3RyICIiCiJBbnbkbmRuaW5nOlxu
IgoiXHQlcyBbLXNdXG4iCgojOiBzcmMva2JkX21vZGUuYzoxOAptc2dpZCAidXNhZ2U6IGtiZF9t
b2RlIFstYXwtdXwta3wtc11cbiIKbXNnc3RyICJhbnbkbmRuaW5nOiBrYmRfbW9kZSBbLWF8LXV8
LWt8LXNdXG4iCgojOiBzcmMva2JkX21vZGUuYzo0MQptc2dpZCAia2JkX21vZGU6IGVycm9yIHJl
YWRpbmcga2V5Ym9hcmQgbW9kZVxuIgptc2dzdHIgImtiZF9tb2RlOiBmZWwgdmlkIGzkc25pbmcg
YXYgdGFuZ2VudGJvcmRzbORnZVxuIgoKIzogc3JjL2tiZF9tb2RlLmM6NDYKbXNnaWQgIlRoZSBr
ZXlib2FyZCBpcyBpbiByYXcgKHNjYW5jb2RlKSBtb2RlXG4iCm1zZ3N0ciAiVGFuZ2VudGJvcmRl
dCDkciBpIHLldHQgKGF2bORzbmluZ3Nrb2RzLSls5GdlXG4iCgojOiBzcmMva2JkX21vZGUuYzo0
OQptc2dpZCAiVGhlIGtleWJvYXJkIGlzIGluIG1lZGl1bXJhdyAoa2V5Y29kZSkgbW9kZVxuIgpt
c2dzdHIgIlRhbmdlbnRib3JkZXQg5HIgaSBoYWx2cuV0dCAodGFuZ2VudGtvZHMtKWzkZ2VcbiIK
CiM6IHNyYy9rYmRfbW9kZS5jOjUyCm1zZ2lkICJUaGUga2V5Ym9hcmQgaXMgaW4gdGhlIGRlZmF1
bHQgKEFTQ0lJKSBtb2RlXG4iCm1zZ3N0ciAiVGFuZ2VudGJvcmRldCDkciBpIHN0YW5kYXJkbORn
ZSAoQVNDSUkpXG4iCgojOiBzcmMva2JkX21vZGUuYzo1NQptc2dpZCAiVGhlIGtleWJvYXJkIGlz
IGluIFVuaWNvZGUgKFVURi04KSBtb2RlXG4iCm1zZ3N0ciAiVGFuZ2VudGJvcmRldCDkciBpIFVu
aWNvZGVs5GdlIChVVEYtOClcbiIKCiM6IHNyYy9rYmRfbW9kZS5jOjU4Cm1zZ2lkICJUaGUga2V5
Ym9hcmQgaXMgaW4gc29tZSB1bmtub3duIG1vZGVcbiIKbXNnc3RyICJUYW5nZW50Ym9yZGV0IORy
IGkgbuVnb3Qgb2vkbnQgbORnZVxuIgoKIzogc3JjL2tiZF9tb2RlLmM6NzYKIywgYy1mb3JtYXQK
bXNnaWQgIiVzOiBlcnJvciBzZXR0aW5nIGtleWJvYXJkIG1vZGVcbiIKbXNnc3RyICIlczogZmVs
IG7kciB0YW5nZW50Ym9yZHNs5GdlIHNhdHRlc1xuIgoKIzogc3JjL2tiZHJhdGUuYzoxMzkgc3Jj
L2tiZHJhdGUuYzoyNzgKIywgYy1mb3JtYXQKbXNnaWQgIlR5cGVtYXRpYyBSYXRlIHNldCB0byAl
LjFmIGNwcyAoZGVsYXkgPSAlZCBtcylcbiIKbXNnc3RyICJVcHByZXBuaW5nc2hhc3RpZ2hldCBz
YXR0IHRpbGwgJS4xZiB0L3MgKGb2cmRy9mpuaW5nID0gJWQgbXMpXG4iCgojOiBzcmMva2JkcmF0
ZS5jOjIyMwptc2dpZCAiVXNhZ2U6IGtiZHJhdGUgWy1WXSBbLXNdIFstciByYXRlXSBbLWQgZGVs
YXldXG4iCm1zZ3N0ciAiQW525G5kbmluZzoga2JkcmF0ZSBbLVZdIFstc10gWy1yIGZyZWt2ZW5z
XSBbLWQgZvZyZHL2am5pbmddXG4iCgojOiBzcmMva2JkcmF0ZS5jOjI1Mwptc2dpZCAiQ2Fubm90
IG9wZW4gL2Rldi9wb3J0Igptc2dzdHIgIkthbiBpbnRlIPZwcG5hIC9kZXYvcG9ydCIKCiM6IHNy
Yy9rZGZvbnRvcC5jOjE5Mwptc2dpZCAiYnVnOiBnZXRmb250IGNhbGxlZCB3aXRoIGNvdW50PDI1
NlxuIgptc2dzdHIgImZlbDogZ2V0Zm9udCBhbnJvcGFkIG1lZCBjb3VudDwyNTZcbiIKCiM6IHNy
Yy9rZGZvbnRvcC5jOjI1MiBzcmMveG1hbGxvYy5jOjE0CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczog
b3V0IG9mIG1lbW9yeVxuIgptc2dzdHIgIiVzOiBtaW5uZXQgc2x1dFxuIgoKIzogc3JjL2tzeW1z
LmM6MTY3MAojLCBjLWZvcm1hdAptc2dpZCAidW5rbm93biBjaGFyc2V0ICVzIC0gaWdub3Jpbmcg
Y2hhcnNldCByZXF1ZXN0XG4iCm1zZ3N0ciAib2vkbmQgdGVja2VudXBwc+R0dG5pbmcgJXMgLSBp
Z25vcmVyYXIgYmVn5HJhbiBvbSB0ZWNrZW51cHBz5HR0bmluZ1xuIgoKIzogc3JjL2tzeW1zLmM6
MTc0MgojLCBjLWZvcm1hdAptc2dpZCAiYXNzdW1pbmcgaXNvLTg4NTktMSAlc1xuIgptc2dzdHIg
ImFudGFyIGlzby04ODU5LTEgJXNcbiIKCiM6IHNyYy9rc3ltcy5jOjE3NDkKIywgYy1mb3JtYXQK
bXNnaWQgImFzc3VtaW5nIGlzby04ODU5LTE1ICVzXG4iCm1zZ3N0ciAiYW50YXIgaXNvLTg4NTkt
MTUgJXNcbiIKCiM6IHNyYy9rc3ltcy5jOjE3NTYKIywgYy1mb3JtYXQKbXNnaWQgImFzc3VtaW5n
IGlzby04ODU5LTIgJXNcbiIKbXNnc3RyICJhbnRhciBpc28tODg1OS0yICVzXG4iCgojOiBzcmMv
a3N5bXMuYzoxNzYzCiMsIGMtZm9ybWF0Cm1zZ2lkICJhc3N1bWluZyBpc28tODg1OS0zICVzXG4i
Cm1zZ3N0ciAiYW50YXIgaXNvLTg4NTktMyAlc1xuIgoKIzogc3JjL2tzeW1zLmM6MTc3MAojLCBj
LWZvcm1hdAptc2dpZCAiYXNzdW1pbmcgaXNvLTg4NTktNCAlc1xuIgptc2dzdHIgImFudGFyIGlz
by04ODU5LTQgJXNcbiIKCiM6IHNyYy9rc3ltcy5jOjE3NzUKIywgYy1mb3JtYXQKbXNnaWQgInVu
a25vd24ga2V5c3ltICclcydcbiIKbXNnc3RyICJva+RuZCB0ZWNrZW5zeW1ib2wgXCIlc1wiXG4i
CgojOiBzcmMva3N5bXMuYzoxODEwCiMsIGMtZm9ybWF0Cm1zZ2lkICJwbHVzIGJlZm9yZSAlcyBp
Z25vcmVkXG4iCm1zZ3N0ciAicGx1cyBm9nJlICVzIGlnbm9yZXJhdFxuIgoKIzogc3JjL2xvYWR1
bmltYXAuYzo2MgojLCBjLWZvcm1hdAptc2dpZCAidXNhZ2U6ICVzIFstbyBtYXAub3JpZ10gW21h
cC1maWxlXVxuIgptc2dzdHIgImFuduRuZG5pbmc6ICVzIFstbyBvcmlnaW5hbHRhYmVsbF0gW3Rh
YmVsbGZpbF1cbiIKCiM6IHNyYy9sb2FkdW5pbWFwLmM6MTUyIHNyYy9sb2FkdW5pbWFwLmM6MTYz
CiMsIGMtZm9ybWF0Cm1zZ2lkICJCYWQgaW5wdXQgbGluZTogJXNcbiIKbXNnc3RyICJGZWxha3Rp
ZyBpbmRhdGFyYWQ6ICVzXG4iCgojOiBzcmMvbG9hZHVuaW1hcC5jOjE3MgojLCBjLWZvcm1hdApt
c2dpZCAiJXM6IEdseXBoIG51bWJlciAoMHgleCkgbGFyZ2VyIHRoYW4gZm9udCBsZW5ndGhcbiIK
bXNnc3RyICIlczogVGVja2VubnVtbWVyICgweCV4KSBzdPZycmUg5G4gdHlwc25pdHRzbORuZ2Rc
biIKCiM6IHNyYy9sb2FkdW5pbWFwLmM6MTc4CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogQmFkIGVu
ZCBvZiByYW5nZSAoMHgleClcbiIKbXNnc3RyICIlczogRmVsYWt0aWd0IHNsdXQgcOUgaW50ZXJ2
YWxsICgweCV4KVxuIgoKIzogc3JjL2xvYWR1bmltYXAuYzoyMDggc3JjL3BzZnh0YWJsZS5jOjE3
NQojLCBjLWZvcm1hdAptc2dpZCAiJXM6IEJhZCBVbmljb2RlIHJhbmdlIGNvcnJlc3BvbmRpbmcg
dG8gZm9udCBwb3NpdGlvbiByYW5nZSAweCV4LTB4JXhcbiIKbXNnc3RyICIlczogRmVsYWt0aWd0
IFVuaWNvZGVpbnRlcnZhbGwgc29tIG1vdHN2YXJhciB0eXBzbml0dHNwb3NpdGlvbnNpbnRlcnZh
bGwgMHgleC0weCV4XG4iCgojOiBzcmMvbG9hZHVuaW1hcC5jOjIxNSBzcmMvcHNmeHRhYmxlLmM6
MTgyCiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogVW5pY29kZSByYW5nZSBVKyV4LVUrJXggbm90IG9m
IHRoZSBzYW1lIGxlbmd0aCBhcyBmb250IHBvc2l0aW9uIHJhbmdlIDB4JXgtMHgleFxuIgptc2dz
dHIgIiVzOiBVbmljb2RlaW50ZXJ2YWxsIFUrJXgtVSsleCDkciBpbnRlIGF2IHNhbW1hIGzkbmdk
IHNvbSB0eXBzbml0dHNwb3NpdGlvbnNpbnRlcnZhbGwgMHgleC0weCV4XG4iCgojOiBzcmMvbG9h
ZHVuaW1hcC5jOjIzNCBzcmMvcHNmeHRhYmxlLmM6MjAzCiMsIGMtZm9ybWF0Cm1zZ2lkICIlczog
dHJhaWxpbmcganVuayAoJXMpIGlnbm9yZWRcbiIKbXNnc3RyICIlczogZWZ0ZXJm9mxqYW5kZSBz
a3LkcCAoJXMpIGlnbm9yZXJhdFxuIgoKIzogc3JjL2xvYWR1bmltYXAuYzoyNTEKIywgYy1mb3Jt
YXQKbXNnaWQgIkxvYWRpbmcgdW5pY29kZSBtYXAgZnJvbSBmaWxlICVzXG4iCm1zZ3N0ciAiTORz
ZXIgaW4gdW5pY29kZXRhYmVsbCBmcuVuIGZpbCAlc1xuIgoKIzogc3JjL2xvYWR1bmltYXAuYzoy
NTcKIywgYy1mb3JtYXQKbXNnaWQgIiVzOiAlczogV2FybmluZzogbGluZSB0b28gbG9uZ1xuIgpt
c2dzdHIgIiVzOiAlczogVmFybmluZzogcmFkZW4g5HIgZvZyIGzlbmdcbiIKCiM6IHNyYy9sb2Fk
dW5pbWFwLmM6MjY3CiMsIGMtZm9ybWF0Cm1zZ2lkICIiCiIlczogbm90IGxvYWRpbmcgZW1wdHkg
dW5pbWFwXG4iCiIoaWYgeW91IGluc2lzdDogdXNlIG9wdGlvbiAtZiB0byBvdmVycmlkZSlcbiIK
bXNnc3RyICIiCiIlczogbORzZXIgaW50ZSBpbiB0b20gdW5pdGFiZWxsXG4iCiIob20gZHUgaW5z
aXN0ZXJhcjogYW525G5kIGZsYWdnYW4gLWYgZvZyIGF0dCDlc2lkb3PkdHRhKVxuIgoKIzogc3Jj
L2xvYWR1bmltYXAuYzoyODgKbXNnaWQgImVudHJ5Igptc2dzdHIgInBvc3QiCgojOiBzcmMvbG9h
ZHVuaW1hcC5jOjI4OAptc2dpZCAiZW50cmllcyIKbXNnc3RyICJwb3N0ZXIiCgojOiBzcmMvbG9h
ZHVuaW1hcC5jOjMxNAojLCBjLWZvcm1hdAptc2dpZCAiU2F2ZWQgdW5pY29kZSBtYXAgb24gYCVz
J1xuIgptc2dzdHIgIlNwYXJhZGUgdW5pY29kZXRhYmVsbCB0aWxsIFwiJXNcIlxuIgoKIzogc3Jj
L2xvYWR1bmltYXAuYzozMzQKbXNnaWQgIkFwcGVuZGVkIFVuaWNvZGUgbWFwXG4iCm1zZ3N0ciAi
TGFkZSB0aWxsIFVuaWNvZGV0YWJlbGxcbiIKCiM6IHNyYy9tYXBzY3JuLmM6NjUKIywgYy1mb3Jt
YXQKbXNnaWQgInVzYWdlOiAlcyBbLXZdIFstbyBtYXAub3JpZ10gbWFwLWZpbGVcbiIKbXNnc3Ry
ICJhbnbkbmRuaW5nOiAlcyBbLXZdIFstbyBvcmlnaW5hbHRhYmVsbF0gdGFiZWxsZmlsXG4iCgoj
OiBzcmMvbWFwc2Nybi5jOjEzMAojLCBjLWZvcm1hdAptc2dpZCAibWFwc2NybjogY2Fubm90IG9w
ZW4gbWFwIGZpbGUgXyVzX1xuIgptc2dzdHIgIm1hcHNjcm46IGthbiBpbnRlIPZwcG5hIHRhYmVs
bGZpbCBfJXNfXG4iCgojOiBzcmMvbWFwc2Nybi5jOjEzNgptc2dpZCAiQ2Fubm90IHN0YXQgbWFw
IGZpbGUiCm1zZ3N0ciAiS2FuIGludGUgdGEgc3RhdHVzIHDlIHRhYmVsbGZpbCIKCiM6IHNyYy9t
YXBzY3JuLmM6MTQxCiMsIGMtZm9ybWF0Cm1zZ2lkICJMb2FkaW5nIGJpbmFyeSBkaXJlY3QtdG8t
Zm9udCBzY3JlZW4gbWFwIGZyb20gZmlsZSAlc1xuIgptc2dzdHIgIkzkc2VyIGluIGJpbuRyIGRp
cmVrdC10aWxsLXR5cHNuaXR0LXNr5HJtdGFiZWxsIGZy5W4gZmlsICVzXG4iCgojOiBzcmMvbWFw
c2Nybi5jOjE0NiBzcmMvbWFwc2Nybi5jOjE1NwojLCBjLWZvcm1hdAptc2dpZCAiRXJyb3IgcmVh
ZGluZyBtYXAgZnJvbSBmaWxlIGAlcydcbiIKbXNnc3RyICJGZWwgdmlkIGzkc25pbmcgYXYgdGFi
ZWxsIGZy5W4gZmlsIFwiJXNcIlxuIgoKIzogc3JjL21hcHNjcm4uYzoxNTIKIywgYy1mb3JtYXQK
bXNnaWQgIkxvYWRpbmcgYmluYXJ5IHVuaWNvZGUgc2NyZWVuIG1hcCBmcm9tIGZpbGUgJXNcbiIK
bXNnc3RyICJM5HNlciBpbiBiaW7kciB1bmljb2RlLXNr5HJtZmlsIGZy5W4gZmlsICVzXG4iCgoj
OiBzcmMvbWFwc2Nybi5jOjE2NAojLCBjLWZvcm1hdAptc2dpZCAiTG9hZGluZyBzeW1ib2xpYyBz
Y3JlZW4gbWFwIGZyb20gZmlsZSAlc1xuIgptc2dzdHIgIkzkc2VyIGluIHN5bWJvbGlzayBza+Ry
bXRhYmVsbCBmcuVuIGZpbCAlc1xuIgoKIzogc3JjL21hcHNjcm4uYzoxNjgKIywgYy1mb3JtYXQK
bXNnaWQgIkVycm9yIHBhcnNpbmcgc3ltYm9saWMgbWFwIGZyb20gYCVzJywgbGluZSAlZFxuIgpt
c2dzdHIgIkZlbCB2aWQgdG9sa25pbmcgYXYgc3ltYm9saXNrIHRhYmVsbCBmcuVuIFwiJXNcIiwg
cmFkICVkXG4iCgojOiBzcmMvbWFwc2Nybi5jOjI3MiBzcmMvbWFwc2Nybi5jOjI3Nwptc2dpZCAi
RXJyb3Igd3JpdGluZyBtYXAgdG8gZmlsZVxuIgptc2dzdHIgIkZlbCB2aWQgc2tyaXZuaW5nIGF2
IHRhYmVsbCB0aWxsIGZpbFxuIgoKIzogc3JjL21hcHNjcm4uYzoyODEKbXNnaWQgIkNhbm5vdCBy
ZWFkIGNvbnNvbGUgbWFwXG4iCm1zZ3N0ciAiS2FuIGludGUgbORzYSBrb25zb2xsdGFiZWxsXG4i
CgojOiBzcmMvbWFwc2Nybi5jOjI4NwojLCBjLWZvcm1hdAptc2dpZCAiU2F2ZWQgc2NyZWVuIG1h
cCBpbiBgJXMnXG4iCm1zZ3N0ciAiU3BhcmFkZSBza+RybXRhYmVsbCBpIFwiJXNcIlxuIgoKIzog
c3JjL3BzZmZvbnRvcC5jOjY2CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogc2hvcnQgdWNzMiB1bmlj
b2RlIHRhYmxlXG4iCm1zZ3N0ciAiJXM6IGtvcnQgdWNzMi11bmljb2RldGFiZWxsXG4iCgojOiBz
cmMvcHNmZm9udG9wLmM6ODcKIywgYy1mb3JtYXQKbXNnaWQgIiVzOiBzaG9ydCB1dGY4IHVuaWNv
ZGUgdGFibGVcbiIKbXNnc3RyICIlczoga29ydCB1dGY4LXVuaWNvZGV0YWJlbGxcbiIKCiM6IHNy
Yy9wc2Zmb250b3AuYzo5MAojLCBjLWZvcm1hdAptc2dpZCAiJXM6IGJhZCB1dGY4XG4iCm1zZ3N0
ciAiJXM6IGZlbGFrdGlnIHV0ZjhcbiIKCiM6IHNyYy9wc2Zmb250b3AuYzo5MwojLCBjLWZvcm1h
dAptc2dpZCAiJXM6IHVua25vd24gdXRmOCBlcnJvclxuIgptc2dzdHIgIiVzOiBva+RudCB1dGY4
LWZlbFxuIgoKIzogc3JjL3BzZmZvbnRvcC5jOjEyNAojLCBjLWZvcm1hdAptc2dpZCAiJXM6IHNo
b3J0IHVuaWNvZGUgdGFibGVcbiIKbXNnc3RyICIlczoga29ydCB1bmljb2RldGFiZWxsXG4iCgoj
OiBzcmMvcHNmZm9udG9wLmM6MjA0CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogRXJyb3IgcmVhZGlu
ZyBpbnB1dCBmb250Igptc2dzdHIgIiVzOiBGZWwgdmlkIGzkc25pbmcgYXYgaW5kYXRhdHlwc25p
dHQiCgojOiBzcmMvcHNmZm9udG9wLmM6MjE4CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogQmFkIGNh
bGwgb2YgcmVhZHBzZmZvbnRcbiIKbXNnc3RyICIlczogRmVsYWt0aWd0IGFucm9wIGF2IHJlYWRw
c2Zmb250XG4iCgojOiBzcmMvcHNmZm9udG9wLmM6MjMzCiMsIGMtZm9ybWF0Cm1zZ2lkICIlczog
VW5zdXBwb3J0ZWQgcHNmIGZpbGUgbW9kZSAoJWQpXG4iCm1zZ3N0ciAiJXM6IHBzZi1maWxs5Gdl
ICglZCkgc3T2ZHMgaW50ZVxuIgoKIzogc3JjL3BzZmZvbnRvcC5jOjI1MQojLCBjLWZvcm1hdApt
c2dpZCAiJXM6IFVuc3VwcG9ydGVkIHBzZiB2ZXJzaW9uICglZClcbiIKbXNnc3RyICIlczogcHNm
LXZlcnNpb24gKCVkKSBzdPZkcyBpbnRlXG4iCgojOiBzcmMvcHNmZm9udG9wLmM6MjY3CiMsIGMt
Zm9ybWF0Cm1zZ2lkICIlczogemVybyBpbnB1dCBmb250IGxlbmd0aD9cbiIKbXNnc3RyICIlczog
bORuZ2QgYXYgaW5kYXRhdHlwc25pdHQg5HIgbm9sbD9cbiIKCiM6IHNyYy9wc2Zmb250b3AuYzoy
NzIKIywgYy1mb3JtYXQKbXNnaWQgIiVzOiB6ZXJvIGlucHV0IGNoYXJhY3RlciBzaXplP1xuIgpt
c2dzdHIgIiVzOiBzdG9ybGVrIGF2IGluZGF0YXRlY2tlbiDkciBub2xsP1xuIgoKIzogc3JjL3Bz
ZmZvbnRvcC5jOjI3OAojLCBjLWZvcm1hdAptc2dpZCAiJXM6IElucHV0IGZpbGU6IGJhZCBpbnB1
dCBsZW5ndGggKCVkKVxuIgptc2dzdHIgIiVzOiBJbmRhdGFmaWw6IG9naWx0aWcgaW5kYXRhbORu
Z2QgKCVkKVxuIgoKIzogc3JjL3BzZmZvbnRvcC5jOjMxMAojLCBjLWZvcm1hdAptc2dpZCAiJXM6
IElucHV0IGZpbGU6IHRyYWlsaW5nIGdhcmJhZ2VcbiIKbXNnc3RyICIlczogSW5kYXRhZmlsOiBl
ZnRlcmb2bGphbmRlIHNrcuRwXG4iCgojOiBzcmMvcHNmZm9udG9wLmM6MzQ4CiMsIGMtZm9ybWF0
Cm1zZ2lkICJhcHBlbmR1bmljb2RlOiBpbGxlZ2FsIHVuaWNvZGUgJXVcbiIKbXNnc3RyICJhcHBl
bmR1bmljb2RlOiBvZ2lsdGlnIHVuaWNvZGUgJXVcbiIKCiM6IHNyYy9wc2Zmb250b3AuYzo0MzQK
bXNnaWQgIkNhbm5vdCB3cml0ZSBmb250IGZpbGUgaGVhZGVyIgptc2dzdHIgIkthbiBpbnRlIHNr
cml2YSB0eXBzbml0dHNmaWxzaHV2dWQiCgojOiBzcmMvcHNmeHRhYmxlLmM6MTA5CiMsIGMtZm9y
bWF0Cm1zZ2lkICIlczogV2FybmluZzogbGluZSB0b28gbG9uZ1xuIgptc2dzdHIgIiVzOiBWYXJu
aW5nOiByYWRlbiDkciBm9nIgbOVuZ1xuIgoKIzogc3JjL3BzZnh0YWJsZS5jOjEyMyBzcmMvcHNm
eHRhYmxlLmM6MTMzCiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogQmFkIGlucHV0IGxpbmU6ICVzXG4i
Cm1zZ3N0ciAiJXM6IEZlbGFrdGlnIGluZGF0YXJhZDogJXNcbiIKCiM6IHNyYy9wc2Z4dGFibGUu
YzoxNDIKIywgYy1mb3JtYXQKbXNnaWQgIiVzOiBHbHlwaCBudW1iZXIgKDB4JWx4KSBwYXN0IGVu
ZCBvZiBmb250XG4iCm1zZ3N0ciAiJXM6IEdseWZudW1tZXIgKDB4JWx4KSBib3J0b20gc2x1dGV0
IGF2IHR5cHNuaXR0ZXRcbiIKCiM6IHNyYy9wc2Z4dGFibGUuYzoxNDcKIywgYy1mb3JtYXQKbXNn
aWQgIiVzOiBCYWQgZW5kIG9mIHJhbmdlICgweCVseClcbiIKbXNnc3RyICIlczogRmVsYWt0aWd0
IHNsdXQgYXYgaW50ZXJ2YWxsICgweCVseClcbiIKCiM6IHNyYy9wc2Z4dGFibGUuYzoxNjYKIywg
Yy1mb3JtYXQKbXNnaWQgIiVzOiBDb3JyZXNwb25kaW5nIHRvIGEgcmFuZ2Ugb2YgZm9udCBwb3Np
dGlvbnMsIHRoZXJlIHNob3VsZCBiZSBhIFVuaWNvZGUgcmFuZ2VcbiIKbXNnc3RyICIlczogVGls
bCBldHQgbW90c3ZhcmFuZGUgaW50ZXJ2YWxsIGF2IHR5cHNuaXR0c3Bvc2l0aW9uZXIgYm9yZGUg
ZGV0IGZpbm5hcyBldHQgVW5pY29kZWludGVydmFsbFxuIgoKIzogc3JjL3BzZnh0YWJsZS5jOjI1
NQojLCBjLWZvcm1hdAptc2dpZCAiIgoiVXNhZ2U6XG4iCiJcdCVzIGluZm9udCBpbnRhYmxlIG91
dGZvbnRcbiIKbXNnc3RyICIiCiJBbnbkbmRuaW5nOlxuIgoiXHQlcyBpbnR5cHNuaXR0IGludGFi
ZWxsIHV0dHlwc25pdHRcbiIKCiM6IHNyYy9wc2Z4dGFibGUuYzoyNjQKIywgYy1mb3JtYXQKbXNn
aWQgIiIKIlVzYWdlOlxuIgoiXHQlcyBpbmZvbnQgW291dHRhYmxlXVxuIgptc2dzdHIgIiIKIkFu
duRuZG5pbmc6XG4iCiJcdCVzIGludHlwc25pdHQgW3V0dGFiZWxsXVxuIgoKIzogc3JjL3BzZnh0
YWJsZS5jOjI3MwojLCBjLWZvcm1hdAptc2dpZCAiIgoiVXNhZ2U6XG4iCiJcdCVzIGluZm9udCBv
dXRmb250XG4iCm1zZ3N0ciAiIgoiQW525G5kbmluZzpcbiIKIlx0JXMgaW50eXBzbml0dCB1dHR5
cHNuaXR0XG4iCgojOiBzcmMvcHNmeHRhYmxlLmM6Mjk4CiMsIGMtZm9ybWF0Cm1zZ2lkICIiCiJV
c2FnZTpcbiIKIlx0JXMgWy1pIGluZm9udF0gWy1vIG91dGZvbnRdIFstaXQgaW50YWJsZV0gWy1v
dCBvdXR0YWJsZV0gWy1udF1cbiIKbXNnc3RyICIiCiJBbnbkbmRuaW5nOlxuIgoiXHQlcyBbLWkg
aW50eXBzbml0dF0gWy1vIHV0dHlwc25pdHRdIFstaXQgaW50YWJlbGxdIFstb3QgdXR0YWJlbGxd
IFstbnRdXG4iCgojOiBzcmMvcHNmeHRhYmxlLmM6MzU4CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczog
QmFkIG1hZ2ljIG51bWJlciBvbiAlc1xuIgptc2dzdHIgIiVzOiBGZWxha3RpZ3QgbWFnaXNrdCBu
dW1tZXIgcOUgJXNcbiIKCiM6IHNyYy9wc2Z4dGFibGUuYzozNzcKIywgYy1mb3JtYXQKbXNnaWQg
IiVzOiBwc2YgZmlsZSB3aXRoIHVua25vd24gbWFnaWNcbiIKbXNnc3RyICIlczogcHNmLWZpbCBt
ZWQgb2vkbmQgbWFnaVxuIgoKIzogc3JjL3BzZnh0YWJsZS5jOjM5MwojLCBjLWZvcm1hdAptc2dp
ZCAiJXM6IGlucHV0IGZvbnQgZG9lcyBub3QgaGF2ZSBhbiBpbmRleFxuIgptc2dzdHIgIiVzOiBp
bmRhdGF0eXBzbml0dGV0IGhhciBpbnRlIG7lZ290IGluZGV4XG4iCgojOiBzcmMvcmVzaXplY29u
cy5jOjE1MwojLCBjLWZvcm1hdAptc2dpZCAicmVzaXplY29uczogY2Fubm90IGZpbmQgdmlkZW9t
b2RlIGZpbGUgJXNcbiIKbXNnc3RyICJyZXNpemVjb25zOiBrYW4gaW50ZSBoaXR0YSB2aWRlb2zk
Z2VzZmlsICVzXG4iCgojOiBzcmMvcmVzaXplY29ucy5jOjE3Mgptc2dpZCAiSW52YWxpZCBudW1i
ZXIgb2YgbGluZXNcbiIKbXNnc3RyICJPZ2lsdGlndCBhbnRhbCByYWRlclxuIgoKIzogc3JjL3Jl
c2l6ZWNvbnMuYzoyMzgKIywgYy1mb3JtYXQKbXNnaWQgIk9sZCBtb2RlOiAlZHglZCAgTmV3IG1v
ZGU6ICVkeCVkXG4iCm1zZ3N0ciAiR2FtbWFsdCBs5GdlOiAlZNclZCAgTnl0dCBs5GdlOiAlZNcl
ZFxuIgoKIzogc3JjL3Jlc2l6ZWNvbnMuYzoyNDAKIywgYy1mb3JtYXQKbXNnaWQgIk9sZCAjc2Nh
bmxpbmVzOiAlZCAgTmV3ICNzY2FubGluZXM6ICVkICBDaGFyYWN0ZXIgaGVpZ2h0OiAlZFxuIgpt
c2dzdHIgIkdhbW1hbHQgYW50YWwgc2thbm5saW5qZXI6ICVkICBOeXR0IGFudGFsIHNrYW5ubGlu
amVyOiAlZCAgVGVja2VuaPZqZDogJWRcbiIKCiM6IHNyYy9yZXNpemVjb25zLmM6MjUxCiMsIGMt
Zm9ybWF0Cm1zZ2lkICJyZXNpemVjb25zOiB0aGUgY29tbWFuZCBgJXMnIGZhaWxlZFxuIgptc2dz
dHIgInJlc2l6ZWNvbnM6IGtvbW1hbmRvdCBcIiVzXCIgbWlzc2x5Y2thZGVzXG4iCgojOiBzcmMv
cmVzaXplY29ucy5jOjMxOQojLCBjLWZvcm1hdAptc2dpZCAicmVzaXplY29uczogZG9uJ3QgZm9y
Z2V0IHRvIGNoYW5nZSBURVJNIChtYXliZSB0byBjb24lZHglZCBvciBsaW51eC0lZHglZClcbiIK
bXNnc3RyICJyZXNpemVjb25zOiBnbPZtIGludGUg5G5kcmEgVEVSTSAoa2Fuc2tlIHRpbGwgY29u
JWR4JWQgZWxsZXIgbGludXgtJWR4JWQpXG4iCgojOiBzcmMvcmVzaXplY29ucy5jOjMzMgptc2dp
ZCAiIgoicmVzaXplY29uczpcbiIKImNhbGwgaXM6ICByZXNpemVjb25zIENPTFN4Uk9XUyAgb3I6
ICByZXNpemVjb25zIENPTFMgUk9XU1xuIgoib3I6IHJlc2l6ZWNvbnMgLWxpbmVzIFJPV1MsIHdp
dGggUk9XUyBvbmUgb2YgMjUsIDI4LCAzMCwgMzQsIDM2LCA0MCwgNDQsIDUwLCA2MFxuIgptc2dz
dHIgIiIKInJlc2l6ZWNvbnM6XG4iCiJhbnJvcDogcmVzaXplY29ucyBLT0xVTU5FUnhSQURFUiAg
ZWxsZXI6IHJlc2l6ZWNvbnMgS09MVU1ORVIgUkFERVJcbiIKImVsbGVyOiByZXNpemVjb25zIC1s
aW5lcyBSQURFUiwgZORyIFJBREVSIORyIGVuIGF2IDI1LCAyOCwgMzAsIDM0LCAzNiwgNDAsIDQ0
LCA1MCwgNjBcbiIKCiM6IHNyYy9yZXNpemVjb25zLmM6MzcwCm1zZ2lkICJyZXNpemVjb25zOiBj
YW5ub3QgZ2V0IEkvTyBwZXJtaXNzaW9ucy5cbiIKbXNnc3RyICJyZXNpemVjb25zOiBrYW4gaW50
ZSBm5SBJL08tcuR0dGlnaGV0ZXIuXG4iCgojOiBzcmMvc2NyZWVuZHVtcC5jOjQ4Cm1zZ2lkICJ1
c2FnZTogc2NyZWVuZHVtcCBbbl1cbiIKbXNnc3RyICJhbnbkbmRuaW5nOiBzY3JlZW5kdW1wIFtu
XVxuIgoKIzogc3JjL3NjcmVlbmR1bXAuYzo2OAojLCBjLWZvcm1hdAptc2dpZCAiRXJyb3IgcmVh
ZGluZyAlc1xuIgptc2dzdHIgIkZlbCB2aWQgbORzbmluZyBhdiAlc1xuIgoKIzogc3JjL3NjcmVl
bmR1bXAuYzoxMDkKIywgYy1mb3JtYXQKbXNnaWQgImNvdWxkbid0IHJlYWQgJXMsIGFuZCBjYW5u
b3QgaW9jdGwgZHVtcFxuIgptc2dzdHIgImt1bmRlIGludGUgbORzYSAlcywgb2NoIGthbiBpbnRl
IGv2cmEgXCJpb2N0bCBkdW1wXCJcbiIKCiMuIHdlIHRyaWVkIHRoaXMganVzdCB0byBiZSBzdXJl
LCBidXQgVElPQ0xJTlVYCiMuIGZ1bmN0aW9uIDAgaGFzIGJlZW4gZGlzYWJsZWQgc2luY2UgMS4x
LjkyCiMuIERvIG5vdCBtZW50aW9uIGBpb2N0bCBkdW1wJyBpbiBlcnJvciBtc2cKIzogc3JjL3Nj
cmVlbmR1bXAuYzoxMTUKIywgYy1mb3JtYXQKbXNnaWQgImNvdWxkbid0IHJlYWQgJXNcbiIKbXNn
c3RyICJrdW5kZSBpbnRlIGzkc2EgJXNcbiIKCiM6IHNyYy9zY3JlZW5kdW1wLmM6MTI0CiMsIGMt
Zm9ybWF0Cm1zZ2lkICJTdHJhbmdlIC4uLiBzY3JlZW4gaXMgYm90aCAlZHglZCBhbmQgJWR4JWQg
Pz9cbiIKbXNnc3RyICJLb25zdGlndCAuLi4gc2vkcm1lbiDkciBi5WRlICVk1yVkIG9jaCAlZNcl
ZD8/XG4iCgojOiBzcmMvc2NyZWVuZHVtcC5jOjE0Mgptc2dpZCAiRXJyb3Igd3JpdGluZyBzY3Jl
ZW5kdW1wXG4iCm1zZ3N0ciAiRmVsIHZpZCBza3Jpdm5pbmcgYXYgc2vkcm1kdW1wXG4iCgojOiBz
cmMvc2V0Zm9udC5jOjczCm1zZ2lkICIiCiJVc2FnZTogc2V0Zm9udCBbd3JpdGUtb3B0aW9uc10g
Wy08Tj5dIFtuZXdmb250Li5dIFstbSBjb25zb2xlbWFwXSBbLXUgdW5pY29kZW1hcF1cbiIKIiAg
d3JpdGUtb3B0aW9ucyAodGFrZSBwbGFjZSBiZWZvcmUgZmlsZSBsb2FkaW5nKTpcbiIKIiAgICAt
byAgPGZpbGVuYW1lPlx0V3JpdGUgY3VycmVudCBmb250IHRvIDxmaWxlbmFtZT5cbiIKIiAgICAt
TyAgPGZpbGVuYW1lPlx0V3JpdGUgY3VycmVudCBmb250IGFuZCB1bmljb2RlIG1hcCB0byA8Zmls
ZW5hbWU+XG4iCiIgICAgLW9tIDxmaWxlbmFtZT5cdFdyaXRlIGN1cnJlbnQgY29uc29sZW1hcCB0
byA8ZmlsZW5hbWU+XG4iCiIgICAgLW91IDxmaWxlbmFtZT5cdFdyaXRlIGN1cnJlbnQgdW5pY29k
ZW1hcCB0byA8ZmlsZW5hbWU+XG4iCiJJZiBubyBuZXdmb250IGFuZCBubyAtW298T3xvbXxvdXxt
fHVdIG9wdGlvbiBpcyBnaXZlbixcbiIKImEgZGVmYXVsdCBmb250IGlzIGxvYWRlZDpcbiIKIiAg
ICBzZXRmb250ICAgICAgICAgICAgIExvYWQgZm9udCBcImRlZmF1bHRbLmd6XVwiXG4iCiIgICAg
c2V0Zm9udCAtPE4+ICAgICAgICBMb2FkIGZvbnQgXCJkZWZhdWx0OHg8Tj5bLmd6XVwiXG4iCiJU
aGUgLTxOPiBvcHRpb24gc2VsZWN0cyBhIGZvbnQgZnJvbSBhIGNvZGVwYWdlIHRoYXQgY29udGFp
bnMgdGhyZWUgZm9udHM6XG4iCiIgICAgc2V0Zm9udCAtezh8MTR8MTZ9IGNvZGVwYWdlLmNwWy5n
el0gICBMb2FkIDh4PE4+IGZvbnQgZnJvbSBjb2RlcGFnZS5jcFxuIgoiRXhwbGljaXRseSAod2l0
aCAtbSBvciAtdSkgb3IgaW1wbGljaXRseSAoaW4gdGhlIGZvbnRmaWxlKSBnaXZlbiBtYXBwaW5n
c1xuIgoid2lsbCBiZSBsb2FkZWQgYW5kLCBpbiB0aGUgY2FzZSBvZiBjb25zb2xlbWFwcywgYWN0
aXZhdGVkLlxuIgoiICAgIC1oPE4+ICAgICAgKG5vIHNwYWNlKSBPdmVycmlkZSBmb250IGhlaWdo
dC5cbiIKIiAgICAtbSA8Zm4+ICAgIExvYWQgY29uc29sZSBzY3JlZW4gbWFwLlxuIgoiICAgIC11
IDxmbj4gICAgTG9hZCBmb250IHVuaWNvZGUgbWFwLlxuIgoiICAgIC1tIG5vbmVcdFN1cHByZXNz
IGxvYWRpbmcgYW5kIGFjdGl2YXRpb24gb2YgYSBzY3JlZW4gbWFwLlxuIgoiICAgIC11IG5vbmVc
dFN1cHByZXNzIGxvYWRpbmcgb2YgYSB1bmljb2RlIG1hcC5cbiIKIiAgICAtdlx0XHRCZSB2ZXJi
b3NlLlxuIgoiICAgIC1WXHRcdFByaW50IHZlcnNpb24gYW5kIGV4aXQuXG4iCiJGaWxlcyBhcmUg
bG9hZGVkIGZyb20gdGhlIGN1cnJlbnQgZGlyZWN0b3J5IG9yIC91c3IvbGliL2tiZC8qLy5cbiIK
bXNnc3RyICIiCiJBbnbkbmRuaW5nOiBzZXRmb250IFtza3JpdmZsYWdnb3JdIFstPE4+XSBbbnl0
dHlwc25pdHQuLl0gWy1tIGtvbnNvbGx0YWJlbGxdIFstdSB1bmljb2RldGFiZWxsXVxuIgoiICBz
a3JpdmZsYWdnb3IgKGjkbmRlciBm9nJlIGZpbGVyIGzkc2VzKTpcbiIKIiAgICAtbyAgPGZpbG5h
bW4+XHRTa3JpdiBudXZhcmFuZGUgdHlwc25pdHQgdGlsbCA8ZmlsbmFtbj5cbiIKIiAgICAtTyAg
PGZpbG5hbW4+XHRTa3JpdiBudXZhcmFuZGUgdHlwc25pdHQgb2NoIHVuaWNvZGV0YWJlbGwgdGls
bCA8ZmlsbmFtbj5cbiIKIiAgICAtb20gPGZpbG5hbW4+XHRTa3JpdiBudXZhcmFuZGUga29uc29s
bHRhYmVsbCB0aWxsIDxmaWxuYW1uPlxuIgoiICAgIC1vdSA8ZmlsbmFtbj5cdFNrcml2IG51dmFy
YW5kZSB1bmljb2RldGFiZWxsIHRpbGwgPGZpbG5hbW4+XG4iCiJPbSBpbmdldCBcIm55dHR5cHNu
aXR0XCIgb2NoIGluZ2VuIC1bb3xPfG9tfG91fG18dV0tZmxhZ2dhIORyIGdpdmVuLFxuIgoibORz
ZXMgZXR0IHN0YW5kYXJkdHlwc25pdHQgaW46XG4iCiIgICAgc2V0Zm9udCAgICAgICAgICAgICBM
5HMgaW4gdHlwc25pdHQgXCJkZWZhdWx0Wy5nel1cIlxuIgoiICAgIHNldGZvbnQgLTxOPiAgICAg
ICAgTORzIGluIHR5cHNuaXR0IFwiZGVmYXVsdDh4PE4+Wy5nel1cIlxuIgoiLTxOPi1mbGFnZ2Fu
IHbkbGplciBldHQgdHlwc25pdHQgZnLlbiBlbiB0ZWNrZW50YWJlbGwgc29tIGlubmVo5WxsZXIg
dHJlIHR5cHNuaXR0OlxuIgoiICAgIHNldGZvbnQgLXs4fDE0fDE2fSBjb2RlcGFnZS5jcFsuZ3pd
ICAgTORzIGluIDjXPE4+LXR5cHNuaXR0IGZy5W4gY29kZXBhZ2UuY3BcbiIKIkV4cGxpY2l0ICht
ZWQgLW0gZWxsZXIgLXUpIGVsbGVyIGltcGxpY2l0IChpIHR5cHNuaXR0c2ZpbGVuKSBnaXZuYSB0
YWJlbGxlclxuIgoia29tbWVyIGzkc2FzIGluIG9jaCwgb20gZGV0IGfkbGxlciBrb25zb2xsdGFi
ZWxsZXIsIGFrdGl2ZXJhcy5cbiIKIiAgICAtaDxOPiAgICAgIChpbmdldCBibGFua3RlY2tlbikg
5XNpZG9z5HR0IHR5cHNuaXR0c2j2amQuXG4iCiIgICAgLW0gPGZuPiAgICBM5HMgaW4ga29uc29s
bHNr5HJtc3RhYmVsbC5cbiIKIiAgICAtdSA8Zm4+ICAgIEzkcyBpbiB1bmljb2RldHlwc25pdHRz
dGFiZWxsLlxuIgoiICAgIC1tIG5vbmVcdEzldCBibGkgYXR0IGzkc2EgaW4gb2NoIGFrdGl2ZXJh
IHNr5HJtdGFiZWxsLlxuIgoiICAgIC11IG5vbmVcdEzldCBibGkgYXR0IGzkc2EgaW4gdW5pY29k
ZXRhYmVsbC5cbiIKIiAgICAtdlx0XHRWYXIgcHJhdHNhbS5cbiIKIiAgICAtVlx0XHRTa3JpdiB1
dCB2ZXJzaW9uIG9jaCBhdnNsdXRhLlxuIgoiRmlsZXIgbORzZXMgaW4gZnLlbiBkZW4gYWt0dWVs
bGEga2F0YWxvZ2VuIGVsbGVyIC91c3IvbGliL2tiZC8qLy5cbiIKCiM6IHNyYy9zZXRmb250LmM6
MTY5Cm1zZ2lkICJzZXRmb250OiB0b28gbWFueSBpbnB1dCBmaWxlc1xuIgptc2dzdHIgInNldGZv
bnQ6IGb2ciBt5W5nYSBpbmRhdGFmaWxlclxuIgoKIzogc3JjL3NldGZvbnQuYzoxNzcKbXNnaWQg
InNldGZvbnQ6IGNhbm5vdCBib3RoIHJlc3RvcmUgZnJvbSBjaGFyYWN0ZXIgUk9NIGFuZCBmcm9t
IGZpbGUuIEZvbnQgdW5jaGFuZ2VkLlxuIgptc2dzdHIgInNldGZvbnQ6IGthbiBpbnRlIGLlZGUg
5XRlcnN05GxsYSBmcuVuIHRlY2tlbi1ST00gb2NoIGZy5W4gZmlsLiBGb250ZW4gb2b2cuRuZHJh
ZC5cbiIKCiM6IHNyYy9zZXRmb250LmM6MjM2CiMsIGMtZm9ybWF0Cm1zZ2lkICJCYWQgY2hhcmFj
dGVyIGhlaWdodCAlZFxuIgptc2dzdHIgIkZlbGFrdGlnIHRlY2tlbmj2amQgJWRcbiIKCiM6IHNy
Yy9zZXRmb250LmM6MjQwCiMsIGMtZm9ybWF0Cm1zZ2lkICJCYWQgY2hhcmFjdGVyIHdpZHRoICVk
XG4iCm1zZ3N0ciAiRmVsYWt0aWcgdGVja2VuYnJlZGQgJWRcbiIKCiM6IHNyYy9zZXRmb250LmM6
MjY1CiMsIGMtZm9ybWF0Cm1zZ2lkICIlczogZm9udCBwb3NpdGlvbiAzMiBpcyBub25ibGFua1xu
Igptc2dzdHIgIiVzOiBUeXBzbml0dHNwb3NpdGlvbiAzMiDkciBpY2tlLWJsYW5rXG4iCgojOiBz
cmMvc2V0Zm9udC5jOjI3MwojLCBjLWZvcm1hdAptc2dpZCAiJXM6IHdpcGVkIGl0XG4iCm1zZ3N0
ciAiJXM6IHJlbnNhZGUgZGV0XG4iCgojOiBzcmMvc2V0Zm9udC5jOjI3NwojLCBjLWZvcm1hdApt
c2dpZCAiJXM6IGJhY2tncm91bmQgd2lsbCBsb29rIGZ1bm55XG4iCm1zZ3N0ciAiJXM6IGJha2dy
dW5kZW4ga29tbWVyIHNlIGtvbnN0aWcgdXRcbiIKCiM6IHNyYy9zZXRmb250LmM6Mjg3CiMsIGMt
Zm9ybWF0Cm1zZ2lkICJMb2FkaW5nICVkLWNoYXIgJWR4JWQgZm9udCBmcm9tIGZpbGUgJXNcbiIK
bXNnc3RyICJM5HNlciBpbiAlZC10ZWNrZW5zICVk1yVkLXR5cHNuaXR0IGZy5W4gZmlsZW4gJXNc
biIKCiM6IHNyYy9zZXRmb250LmM6MjkwCiMsIGMtZm9ybWF0Cm1zZ2lkICJMb2FkaW5nICVkLWNo
YXIgJWR4JWQgZm9udFxuIgptc2dzdHIgIkzkc2VyIGluICVkLXRlY2tlbnMgJWTXJWQtdHlwc25p
dHRcbiIKCiM6IHNyYy9zZXRmb250LmM6MjkzCiMsIGMtZm9ybWF0Cm1zZ2lkICJMb2FkaW5nICVk
LWNoYXIgJWR4JWQgKCVkKSBmb250IGZyb20gZmlsZSAlc1xuIgptc2dzdHIgIkzkc2VyIGluICVk
LXRlY2tlbnMgJWTXJWQtdHlwc25pdHQgKCVkKSBmcuVuIGZpbGVuICVzXG4iCgojOiBzcmMvc2V0
Zm9udC5jOjI5NgojLCBjLWZvcm1hdAptc2dpZCAiTG9hZGluZyAlZC1jaGFyICVkeCVkICglZCkg
Zm9udFxuIgptc2dzdHIgIkzkc2VyIGluICVkLXRlY2tlbnMgJWTXJWQtdHlwc25pdHQgKCVkKVxu
IgoKIzogc3JjL3NldGZvbnQuYzozMzYKIywgYy1mb3JtYXQKbXNnaWQgIiVzOiBidWcgaW4gZG9f
bG9hZHRhYmxlXG4iCm1zZ3N0ciAiJXM6IGZlbCBpIGRvX2xvYWR0YWJsZVxuIgoKIzogc3JjL3Nl
dGZvbnQuYzozNDIKbXNnaWQgIkxvYWRpbmcgVW5pY29kZSBtYXBwaW5nIHRhYmxlLi4uXG4iCm1z
Z3N0ciAiTORzZXIgaW4gVW5pY29kZS1rb252ZXJ0ZXJpbmdzc3RhYmVsbC4uLlxuIgoKIzogc3Jj
L3NldGZvbnQuYzozNzggc3JjL3NldGZvbnQuYzo0NjIKIywgYy1mb3JtYXQKbXNnaWQgIkNhbm5v
dCBvcGVuIGZvbnQgZmlsZSAlc1xuIgptc2dzdHIgIkthbiBpbnRlIPZwcG5hIHR5cHNuaXR0c2Zp
bGVuICVzXG4iCgojOiBzcmMvc2V0Zm9udC5jOjM4OQojLCBjLWZvcm1hdAptc2dpZCAiV2hlbiBs
b2FkaW5nIHNldmVyYWwgZm9udHMsIGFsbCBtdXN0IGJlIHBzZiBmb250cyAtICVzIGlzbid0XG4i
Cm1zZ3N0ciAiTuRyIGZsZXJhIHR5cHNuaXR0IGzkc2VzIGluIG3lc3RlIGFsbGEgdmFyYSBwc2Yt
dHlwc25pdHQgLSAlcyDkciBpbnRlIGRldFxuIgoKIzogc3JjL3NldGZvbnQuYzozOTcKIywgYy1m
b3JtYXQKbXNnaWQgIlJlYWQgJWQtY2hhciAlZHglZCBmb250IGZyb20gZmlsZSAlc1xuIgptc2dz
dHIgIkzkc3RlICVkLXRlY2tlbnMgJWTXJWQtdHlwc25pdHQgZnLlbiBmaWxlbiAlc1xuIgoKIzog
c3JjL3NldGZvbnQuYzo0MDMKbXNnaWQgIldoZW4gbG9hZGluZyBzZXZlcmFsIGZvbnRzLCBhbGwg
bXVzdCBoYXZlIHRoZSBzYW1lIGhlaWdodFxuIgptc2dzdHIgIk7kciBmbGVyYSB0eXBzbml0dCBs
5HNlcyBpbiBt5XN0ZSBhbGxhIGhhIHNhbW1hIGj2amRcbiIKCiM6IHNyYy9zZXRmb250LmM6NDEw
Cm1zZ2lkICJXaGVuIGxvYWRpbmcgc2V2ZXJhbCBmb250cywgYWxsIG11c3QgaGF2ZSB0aGUgc2Ft
ZSB3aWR0aFxuIgptc2dzdHIgIk7kciBmbGVyYSB0eXBzbml0dCBs5HNlcyBpbiBt5XN0ZSBhbGxh
IGhhIHNhbW1hIGJyZWRkXG4iCgojOiBzcmMvc2V0Zm9udC5jOjQ0OQptc2dpZCAiQ2Fubm90IGZp
bmQgZGVmYXVsdCBmb250XG4iCm1zZ3N0ciAiSGl0dGFyIGludGUgc3RhbmRhcmR0eXBzbml0dGV0
XG4iCgojOiBzcmMvc2V0Zm9udC5jOjQ1NgojLCBjLWZvcm1hdAptc2dpZCAiQ2Fubm90IGZpbmQg
JXMgZm9udFxuIgptc2dzdHIgIkhpdHRhciBpbnRlIHR5cHNuaXR0ZXQgJXNcbiIKCiM6IHNyYy9z
ZXRmb250LmM6NDY4CiMsIGMtZm9ybWF0Cm1zZ2lkICJSZWFkaW5nIGZvbnQgZmlsZSAlc1xuIgpt
c2dzdHIgIkzkc2VyIHR5cHNuaXR0c2ZpbGVuICVzXG4iCgojOiBzcmMvc2V0Zm9udC5jOjUwNgpt
c2dpZCAiTm8gZmluYWwgbmV3bGluZSBpbiBjb21iaW5lIGZpbGVcbiIKbXNnc3RyICJJbmdldCBz
bHV0Z2lsdGlndCBueXJhZHN0ZWNrZW4gaSBrb21iaW5hdGlvbnNmaWxlblxuIgoKIzogc3JjL3Nl
dGZvbnQuYzo1MTIKbXNnaWQgIlRvbyBtYW55IGZpbGVzIHRvIGNvbWJpbmVcbiIKbXNnc3RyICJG
9nIgbeVuZ2EgZmlsZXIgYXR0IGtvbWJpbmVyYVxuIgoKIy4gcmVzdG9yZWZvbnQgLXcgd3JpdGVz
IGEgU1ZHQSBmb250IHRvIGZpbGUKIy4gcmVzdG9yZWZvbnQgLXIgcmVzdG9yZXMgaXQKIy4gVGhl
c2UgZm9udHMgaGF2ZSBzaXplIDMyNzY4LCBmb3IgdHdvIDUxMi1jaGFyIGZvbnRzLgojLiBJbiBm
YWN0LCB3aGVuIEJST0tFTl9HUkFQSElDU19QUk9HUkFNUyBpcyBkZWZpbmVkLAojLiBhbmQgaXQg
YWx3YXlzIGlzLCB0aGVyZSBpcyBubyBkZWZhdWx0IGZvbnQgdGhhdCBpcyBzYXZlZCwKIy4gc28g
cHJvYmFibHkgdGhlIHNlY29uZCBoYWxmIGlzIGFsd2F5cyBnYXJiYWdlLgojOiBzcmMvc2V0Zm9u
dC5jOjUzNgptc2dpZCAiSG1tIC0gYSBmb250IGZyb20gcmVzdG9yZWZvbnQ/IFVzaW5nIHRoZSBm
aXJzdCBoYWxmLlxuIgptc2dzdHIgIkhtbSAtIGV0dCB0eXBzbml0dCBmcuVuIHJlc3RvcmVmb250
PyBBbnbkbmRlciBm9nJzdGEgaGFsdmFuLlxuIgoKIzogc3JjL3NldGZvbnQuYzo1NTMKbXNnaWQg
IkJhZCBpbnB1dCBmaWxlIHNpemVcbiIKbXNnc3RyICJGZWxha3RpZyBzdG9ybGVrIHDlIGluZGF0
YWZpbGVuXG4iCgojOiBzcmMvc2V0Zm9udC5jOjU3NAptc2dpZCAiIgoiVGhpcyBmaWxlIGNvbnRh
aW5zIDMgZm9udHM6IDh4OCwgOHgxNCBhbmQgOHgxNi4gUGxlYXNlIGluZGljYXRlXG4iCiJ1c2lu
ZyBhbiBvcHRpb24gLTggb3IgLTE0IG9yIC0xNiB3aGljaCBvbmUgeW91IHdhbnQgbG9hZGVkLlxu
Igptc2dzdHIgIiIKIkRlbiBo5HIgZmlsZW4gaW5uZWjlbGxlciAzIHR5cHNuaXR0OiA41zgsIDjX
MTQgb2NoIDjXMTYuIFbkbGogdmlsa2V0XG4iCiJkdSB2aWxsIGzkc2EgaW4gbWVkIG7lZ29uIGF2
IGZsYWdnb3JuYSAtOCwgLTE0IG9jaCAtMTYuXG4iCgojOiBzcmMvc2V0Zm9udC5jOjU4OAojLCBj
LWZvcm1hdAptc2dpZCAiWW91IGFza2VkIGZvciBmb250IHNpemUgJWQsIGJ1dCBvbmx5IDgsIDE0
LCAxNiBhcmUgcG9zc2libGUgaGVyZS5cbiIKbXNnc3RyICJEdSBiYWQgb20gdHlwc25pdHRzc3Rv
cmxla2VuICVkLCBtZW4gYmFyYSA4LCAxNCBvY2ggMTYg5HIgbfZqbGlnYSBo5HIuXG4iCgojOiBz
cmMvc2V0Zm9udC5jOjYzMwptc2dpZCAiRm91bmQgbm90aGluZyB0byBzYXZlXG4iCm1zZ3N0ciAi
SGl0dGFkZSBpbmdldCBhdHQgc3BhcmFcbiIKCiM6IHNyYy9zZXRmb250LmM6NjM3Cm1zZ2lkICJD
YW5ub3Qgd3JpdGUgZm9udCBmaWxlIgptc2dzdHIgIkthbiBpbnRlIHNrcml2YSB0aWxsIHR5cHNu
aXR0c2ZpbGVuIgoKIzogc3JjL3NldGZvbnQuYzo2NDIKIywgYy1mb3JtYXQKbXNnaWQgIlNhdmVk
ICVkLWNoYXIgJWR4JWQgZm9udCBmaWxlIG9uICVzXG4iCm1zZ3N0ciAiU3BhcmFkZSAlZC10ZWNr
ZW5zICVk1yVkLXR5cHNuaXR0c2ZpbCB0aWxsICVzXG4iCgojOiBzcmMvc2V0a2V5Y29kZXMuYzoy
MQptc2dpZCAiIgoidXNhZ2U6IHNldGtleWNvZGUgc2NhbmNvZGUga2V5Y29kZSAuLi5cbiIKIiAo
d2hlcmUgc2NhbmNvZGUgaXMgZWl0aGVyIHh4IG9yIGUweHgsIGdpdmVuIGluIGhleGFkZWNpbWFs
LFxuIgoiICBhbmQga2V5Y29kZSBpcyBnaXZlbiBpbiBkZWNpbWFsKVxuIgptc2dzdHIgIiIKImFu
duRuZG5pbmc6IHNldGtleWNvZGUgYXZs5HNuaW5nc2tvZCB0YW5nZW50a29kIC4uLlxuIgoiIChk
5HIgYXZs5HNuaW5nc2tvZCDkciBhbnRpbmdlbiB4eCBlbGxlciBlMHh4IGFuZ2l2ZXQgaGV4YWRl
Y2ltYWx0LFxuIgoiICBvY2ggdGFuZ2VudGtvZCDkciBhbmdpdmV0IGRlY2ltYWx0KVxuIgoKIzog
c3JjL3NldGtleWNvZGVzLmM6NDMKbXNnaWQgImV2ZW4gbnVtYmVyIG9mIGFyZ3VtZW50cyBleHBl
Y3RlZCIKbXNnc3RyICJq5G1udCBhbnRhbCBhcmd1bWVudCBm9nJ25G50YWRlcyIKCiM6IHNyYy9z
ZXRrZXljb2Rlcy5jOjUwCm1zZ2lkICJlcnJvciByZWFkaW5nIHNjYW5jb2RlIgptc2dzdHIgImZl
bCB2aWQgbORzbmluZyBhdiBhdmzkc25pbmdza29kIgoKIzogc3JjL3NldGtleWNvZGVzLmM6NTYK
bXNnaWQgImNvZGUgb3V0c2lkZSBib3VuZHMiCm1zZ3N0ciAia29kIHV0YW5m9nIgZ3LkbnNlcm5h
IgoKIzogc3JjL3NldGtleWNvZGVzLmM6NTkKIywgYy1mb3JtYXQKbXNnaWQgImZhaWxlZCB0byBz
ZXQgc2NhbmNvZGUgJXggdG8ga2V5Y29kZSAlZFxuIgptc2dzdHIgImt1bmRlIGludGUgc+R0dGEg
YXZs5HNuaW5nc2tvZGVuICV4IHRpbGwgdGFuZ2VudGtvZGVuICVkXG4iCgojOiBzcmMvc2V0bGVk
cy5jOjI1CiMsIGMtZm9ybWF0Cm1zZ2lkICIiCiJVc2FnZTpcbiIKIlx0c2V0bGVkcyBbLXZdIFst
TF0gWy1EXSBbLUZdIFtbK3wtXVsgbnVtIHwgY2FwcyB8IHNjcm9sbCAlc11dXG4iCiJUaHVzLFxu
IgoiXHRzZXRsZWRzICtjYXBzIC1udW1cbiIKIndpbGwgc2V0IENhcHNMb2NrLCBjbGVhciBOdW1M
b2NrIGFuZCBsZWF2ZSBTY3JvbGxMb2NrIHVuY2hhbmdlZC5cbiIKIlRoZSBzZXR0aW5ncyBiZWZv
cmUgYW5kIGFmdGVyIHRoZSBjaGFuZ2UgKGlmIGFueSkgYXJlIHJlcG9ydGVkXG4iCiJ3aGVuIHRo
ZSAtdiBvcHRpb24gaXMgZ2l2ZW4gb3Igd2hlbiBubyBjaGFuZ2UgaXMgcmVxdWVzdGVkLlxuIgoi
Tm9ybWFsbHksIHNldGxlZHMgaW5mbHVlbmNlcyB0aGUgdnQgZmxhZyBzZXR0aW5nc1xuIgoiKGFu
ZCB0aGVzZSBhcmUgdXN1YWxseSByZWZsZWN0ZWQgaW4gdGhlIGxlZHMpLlxuIgoiV2l0aCAtTCwg
c2V0bGVkcyBvbmx5IHNldHMgdGhlIGxlZHMsIGFuZCBsZWF2ZXMgdGhlIGZsYWdzIGFsb25lLlxu
IgoiV2l0aCAtRCwgc2V0bGVkcyBzZXRzIGJvdGggdGhlIGZsYWdzIGFuZCB0aGUgZGVmYXVsdCBm
bGFncywgc29cbiIKInRoYXQgYSBzdWJzZXF1ZW50IHJlc2V0IHdpbGwgbm90IGNoYW5nZSB0aGUg
ZmxhZ3MuXG4iCm1zZ3N0ciAiIgoiQW525G5kbmluZzpcbiIKIlx0c2V0bGVkcyBbLXZdIFstTF0g
Wy1EXSBbLUZdIFtbK3wtXVsgbnVtIHwgY2FwcyB8IHNjcm9sbCAlc11dXG4iCiJEdnMsXG4iCiJc
dHNldGxlZHMgK2NhcHMgLW51bVxuIgoia29tbWVyIHPkdHRhIGNhcHNsb2NrLCBzdORuZ2EgYXYg
bnVtbG9jayBvY2ggbORtbmEgc2Nyb2xsb2NrIG9m9nLkbmRyYWQuXG4iCiJJbnN05GxsbmluZ2Fy
bmEgZvZyZSBvY2ggZWZ0ZXIg5G5kcmluZyAob20gbuVnb24pIHJhcHBvcnRlcmFzIG7kclxuIgoi
LXYtZmxhZ2dhbiDkciBnaXZlbiBlbGxlciBu5HIgaW5nYSDkbmRyaW5nYXIgYmVn5HJzLlxuIgoi
Tm9ybWFsdCBw5XZlcmthciBzZXRsZWRzIHZ0LWZsYWdnaW5zdORsbG5pbmdhcm5hXG4iCiIob2No
IGRldHRhIHZpc2FzIG5vcm1hbHQgbWVkIGRpb2Rlcm5hKS5cbiIKIk1lZCAtTCBz5HR0ZXIgc2V0
bGVkcyBkaW9kZXJuYSBvY2ggcOV2ZXJrYXIgaW50ZSBmbGFnZ29ybmEuXG4iCiJNZWQgLUQgc+R0
dGVyIGLlZGUgZmxhZ2dvcm5hIG9jaCBzdGFuZGFyZGZsYWdnb3JuYSBz5SBhdHQgc2VuYXJlXG4i
CiJub2xsc3TkbGxuaW5nYXIgaW50ZSBrb21tZXIg5G5kcmEgZmxhZ2dvcm5hLlxuIgoKIzogc3Jj
L3NldGxlZHMuYzo0Nwptc2dpZCAib24gIgptc2dzdHIgInDlIgoKIzogc3JjL3NldGxlZHMuYzo0
Nwptc2dpZCAib2ZmIgptc2dzdHIgImF2IgoKIzogc3JjL3NldGxlZHMuYzo5MAptc2dpZCAiRXJy
b3IgcmVhZGluZyBjdXJyZW50IGxlZCBzZXR0aW5nLiBNYXliZSBzdGRpbiBpcyBub3QgYSBWVD9c
biIKbXNnc3RyICJGZWwgdmlkIGzkc25pbmcgYXYgbnV2YXJhbmRlIGluc3TkbGxuaW5nLiBTdGFu
ZGFyZCBpbiBrYW5za2UgaW50ZSDkciBlbiBWVD9cbiIKCiM6IHNyYy9zZXRsZWRzLmM6MTA5Cm1z
Z2lkICJFcnJvciByZWFkaW5nIGN1cnJlbnQgZmxhZ3Mgc2V0dGluZy4gTWF5YmUgeW91IGFyZSBu
b3Qgb24gdGhlIGNvbnNvbGU/XG4iCm1zZ3N0ciAiRmVsIHZpZCBs5HNuaW5nIGF2IG51dmFyYW5k
ZSBmbGFnZ2luc3TkbGxuaW5nLiBEdSBrYW5za2UgaW50ZSDkciBw5SBrb25zb2xsZW4/XG4iCgoj
OiBzcmMvc2V0bGVkcy5jOjEyMyBzcmMvc2V0bGVkcy5jOjEzOAptc2dpZCAiRXJyb3IgcmVhZGlu
ZyBjdXJyZW50IGxlZCBzZXR0aW5nIGZyb20gL2Rldi9rYmQuXG4iCm1zZ3N0ciAiRmVsIHZpZCBs
5HNuaW5nIGF2IG51dmFyYW5kZSBkaW9kaW5zdORsbG5pbmcgZnLlbiAvZGV2L2tiZC5cbiIKCiM6
IHNyYy9zZXRsZWRzLmM6MTI3Cm1zZ2lkICJLSU9DR0xFRCB1bmF2YWlsYWJsZT9cbiIKbXNnc3Ry
ICJLSU9DR0xFRCBpbnRlIHRpbGxn5G5nbGlnP1xuIgoKIzogc3JjL3NldGxlZHMuYzoxNDIKbXNn
aWQgIktJT0NTTEVEIHVuYXZhaWxhYmxlP1xuIgptc2dzdHIgIktJT0NTTEVEIGludGUgdGlsbGfk
bmdsaWc/XG4iCgojOiBzcmMvc2V0bGVkcy5jOjE2OQptc2dpZCAiRXJyb3Igb3BlbmluZyAvZGV2
L2tiZC5cbiIKbXNnc3RyICJGZWwgdmlkIPZwcG5hbmRlIGF2IC9kZXYva2JkLlxuIgoKIzogc3Jj
L3NldGxlZHMuYzoyMDEKbXNnaWQgIkVycm9yIHJlc2V0dGluZyBsZWRtb2RlXG4iCm1zZ3N0ciAi
RmVsIHZpZCBub2xsc3TkbGxuaW5nIGF2IGRpb2Rs5GdlXG4iCgojOiBzcmMvc2V0bGVkcy5jOjIx
MAptc2dpZCAiQ3VycmVudCBkZWZhdWx0IGZsYWdzOiAgIgptc2dzdHIgIk51dmFyYW5kZSBzdGFu
ZGFyZGZsYWdnb3I6ICAiCgojOiBzcmMvc2V0bGVkcy5jOjIxNAptc2dpZCAiQ3VycmVudCBmbGFn
czogICAgICAgICAgIgptc2dzdHIgIk51dmFyYW5kZSBmbGFnZ29yOiAgICAgICAgICAiCgojOiBz
cmMvc2V0bGVkcy5jOjIxOAptc2dpZCAiQ3VycmVudCBsZWRzOiAgICAgICAgICAgIgptc2dzdHIg
Ik51dmFyYW5kZSBkaW9kZXI6ICAgICAgICAgICAiCgojOiBzcmMvc2V0bGVkcy5jOjI1NCBzcmMv
c2V0bWV0YW1vZGUuYzo5NAojLCBjLWZvcm1hdAptc2dpZCAidW5yZWNvZ25pemVkIGFyZ3VtZW50
OiBfJXNfXG5cbiIKbXNnc3RyICJva+RudCBhcmd1bWVudDogXyVzX1xuXG4iCgojOiBzcmMvc2V0
bGVkcy5jOjI2Mwptc2dpZCAiT2xkIGRlZmF1bHQgZmxhZ3M6ICAgICIKbXNnc3RyICJHYW1sYSBz
dGFuZGFyZGZsYWdnb3I6ICAgICIKCiM6IHNyYy9zZXRsZWRzLmM6MjY1Cm1zZ2lkICJOZXcgZGVm
YXVsdCBmbGFnczogICAgIgptc2dzdHIgIk55YSBzdGFuZGFyZGZsYWdnb3I6ICAgICAgIgoKIzog
c3JjL3NldGxlZHMuYzoyNzIKbXNnaWQgIk9sZCBmbGFnczogICAgICAgICAgICAiCm1zZ3N0ciAi
R2FtbGEgZmxhZ2dvcjogICAgICAgICAgICAiCgojOiBzcmMvc2V0bGVkcy5jOjI3NAptc2dpZCAi
TmV3IGZsYWdzOiAgICAgICAgICAgICIKbXNnc3RyICJOeWEgZmxhZ2dvcjogICAgICAgICAgICAg
ICIKCiM6IHNyYy9zZXRsZWRzLmM6Mjg4IHNyYy9zZXRsZWRzLmM6Mjk3Cm1zZ2lkICJPbGQgbGVk
czogICAgICAgICAgICAgIgptc2dzdHIgIkdhbWxhIGRpb2RlcjogICAgICAgICAgICAgIgoKIzog
c3JjL3NldGxlZHMuYzoyOTAgc3JjL3NldGxlZHMuYzoyOTkKbXNnaWQgIk5ldyBsZWRzOiAgICAg
ICAgICAgICAiCm1zZ3N0ciAiTnlhIGRpb2RlcjogICAgICAgICAgICAgICAiCgojOiBzcmMvc2V0
bWV0YW1vZGUuYzoyMAptc2dpZCAiIgoiVXNhZ2U6XG4iCiJcdHNldG1ldGFtb2RlIFsgbWV0YWJp
dCB8IG1ldGEgfCBiaXQgfCBlc2NwcmVmaXggfCBlc2MgfCBwcmVmaXggXVxuIgoiRWFjaCB2dCBo
YXMgaGlzIG93biBjb3B5IG9mIHRoaXMgYml0LiBVc2VcbiIKIlx0c2V0bWV0YW1vZGUgW2FyZ10g
PCAvZGV2L3R0eW5cbiIKInRvIGNoYW5nZSB0aGUgc2V0dGluZ3Mgb2YgYW5vdGhlciB2dC5cbiIK
IlRoZSBzZXR0aW5nIGJlZm9yZSBhbmQgYWZ0ZXIgdGhlIGNoYW5nZSBhcmUgcmVwb3J0ZWQuXG4i
Cm1zZ3N0ciAiIgoiQW525G5kbmluZzpcbiIKIlx0c2V0bWV0YW1vZGUgWyBtZXRhYml0IHwgbWV0
YSB8IGJpdCB8IGVzY3ByZWZpeCB8IGVzYyB8IHByZWZpeCBdXG4iCiJWYXJqZSB2dCBoYXIgc2lu
IGVnZW4ga29waWEgYXYgZGVuIGjkciBiaXRlbi4gQW525G5kXG4iCiJcdHNldG1ldGFtb2RlIFth
cmddIDwgL2Rldi90dHluXG4iCiJm9nIgYXR0IORuZHJhIGluc3TkbGxuaW5nZW4gZvZyIGVuIGFu
bmFuIHZ0LlxuIgoiSW5zdORsbG5pbmdlbiBm9nJlIG9jaCBlZnRlciBm9nLkbmRyaW5nZW4gcmFw
cG9ydGVyYXMuXG4iCgojOiBzcmMvc2V0bWV0YW1vZGUuYzozNgptc2dpZCAiTWV0YSBrZXkgc2V0
cyBoaWdoIG9yZGVyIGJpdFxuIgptc2dzdHIgIk1ldGF0YW5nZW50ZW4gc+R0dGVyIGj2Z3N0YSBi
aXRlblxuIgoKIzogc3JjL3NldG1ldGFtb2RlLmM6MzkKbXNnaWQgIk1ldGEga2V5IGdpdmVzIEVz
YyBwcmVmaXhcbiIKbXNnc3RyICJNZXRhdGFuZ2VudGVuIGdlciBlc2MtcHJlZml4XG4iCgojOiBz
cmMvc2V0bWV0YW1vZGUuYzo0Mgptc2dpZCAiU3RyYW5nZSBtb2RlIGZvciBNZXRhIGtleT9cbiIK
bXNnc3RyICJLb25zdGlndCBs5GdlIGb2ciBNZXRhdGFuZ2VudGVuP1xuIgoKIzogc3JjL3NldG1l
dGFtb2RlLmM6NzgKbXNnaWQgIkVycm9yIHJlYWRpbmcgY3VycmVudCBzZXR0aW5nLiBNYXliZSBz
dGRpbiBpcyBub3QgYSBWVD9cbiIKbXNnc3RyICJGZWwgdmlkIGzkc25pbmcgYXYgbnV2YXJhbmRl
IGluc3TkbGxuaW5nLiBTdGFuZGFyZCBpbiBrYW5za2UgaW50ZSDkciBlbiBWVD9cbiIKCiM6IHNy
Yy9zZXRtZXRhbW9kZS5jOjk4Cm1zZ2lkICJvbGQgc3RhdGU6ICAgICIKbXNnc3RyICJnYW1tYWx0
IHRpbGxzdOVuZDogICAgIgoKIzogc3JjL3NldG1ldGFtb2RlLmM6MTA0Cm1zZ2lkICJuZXcgc3Rh
dGU6ICAgICIKbXNnc3RyICJueXR0IHRpbGxzdOVuZDogICAgICAgIgoKIzogc3JjL3NldHZlc2Fi
bGFuay5jOjIxCiMsIGMtZm9ybWF0Cm1zZ2lkICJ1c2FnZTogJXNcbiIKbXNnc3RyICJhbnbkbmRu
aW5nOiAlc1xuIgoKIzogc3JjL3Nob3dmb250LmM6MzAKbXNnaWQgImZhaWxlZCB0byByZXN0b3Jl
IG9yaWdpbmFsIHRyYW5zbGF0aW9uIHRhYmxlXG4iCm1zZ3N0ciAibWlzc2x5Y2thZGVzIG1lZCBh
dHQg5XRlcnN05GxsYSBvcmlnaW5hbPZ2ZXJz5HR0bmluZ3N0YWJlbGxlblxuIgoKIzogc3JjL3No
b3dmb250LmM6MzUKbXNnaWQgImZhaWxlZCB0byByZXN0b3JlIG9yaWdpbmFsIHVuaW1hcFxuIgpt
c2dzdHIgIm1pc3NseWNrYWRlcyBtZWQgYXR0IOV0ZXJzdORsbGEgb3JpZ2luYWx1bml0YWJlbGxc
biIKCiM6IHNyYy9zaG93Zm9udC5jOjUzCm1zZ2lkICJjYW5ub3QgY2hhbmdlIHRyYW5zbGF0aW9u
IHRhYmxlXG4iCm1zZ3N0ciAia2FuIGludGUg5G5kcmEg9nZlcnPkdHRuaW5nc3RhYmVsbGVuXG4i
CgojOiBzcmMvc2hvd2ZvbnQuYzo2MAojLCBjLWZvcm1hdAptc2dpZCAiJXM6IG91dCBvZiBtZW1v
cnk/XG4iCm1zZ3N0ciAiJXM6IHNsdXQgcOUgbWlubmU/XG4iCgojOiBzcmMvc2hvd2ZvbnQuYzox
MDEKbXNnaWQgIiIKInVzYWdlOiBzaG93Zm9udCBbLXZ8LVZdXG4iCiIocHJvYmFibHkgYWZ0ZXIg
bG9hZGluZyBhIGZvbnQgd2l0aCBgc2V0Zm9udCBmb250JylcbiIKbXNnc3RyICIiCiJhbnbkbmRu
aW5nOiBzaG93Zm9udCBbLXZ8LVZdXG4iCiIoZvZybW9kbGlnZW4gZWZ0ZXIgYXR0IGhhIGzkc3Qg
aW4gZXR0IHR5cHNuaXR0IG1lZCBcInNldGZvbnQgdHlwc25pdHRcIilcbiIKCiM6IHNyYy9zaG93
a2V5LmM6NDIKbXNnaWQgIj9VTktOT1dOPyIKbXNnc3RyICI/T0vETlQ/IgoKIzogc3JjL3Nob3dr
ZXkuYzo0NAojLCBjLWZvcm1hdAptc2dpZCAia2IgbW9kZSB3YXMgJXNcbiIKbXNnc3RyICJ0Z2It
bORnZSB2YXIgJXNcbiIKCiM6IHNyYy9zaG93a2V5LmM6NDYKbXNnaWQgIiIKIlsgaWYgeW91IGFy
ZSB0cnlpbmcgdGhpcyB1bmRlciBYLCBpdCBtaWdodCBub3Qgd29ya1xuIgoic2luY2UgdGhlIFgg
c2VydmVyIGlzIGFsc28gcmVhZGluZyAvZGV2L2NvbnNvbGUgXVxuIgptc2dzdHIgIiIKIlsgb20g
ZHUgZ/ZyIGRldCBo5HIgaSBYIGthbnNrZSBkZXQgaW50ZSBmdW5nZXJhclxuIgoiZWZ0ZXJzb20g
WC1zZXJ2ZXJuIG9ja3PlIGzkc2VyIC9kZXYvY29uc29sZSBdXG4iCgojOiBzcmMvc2hvd2tleS5j
OjY1CiMsIGMtZm9ybWF0Cm1zZ2lkICJjYXVnaHQgc2lnbmFsICVkLCBjbGVhbmluZyB1cC4uLlxu
Igptc2dzdHIgImZpY2sgc2lnbmFsZW4gJWQsIHN05GRhciB1cHAuLi5cbiIKCiM6IHNyYy9zaG93
a2V5LmM6NzkKIywgYy1mb3JtYXQKbXNnaWQgIiIKInNob3drZXkgdmVyc2lvbiAlc1xuIgoiXG4i
CiJ1c2FnZTogc2hvd2tleSBbb3B0aW9ucy4uLl1cbiIKIlxuIgoidmFsaWQgb3B0aW9ucyBhcmU6
XG4iCiJcbiIKIlx0LWggLS1oZWxwXHRkaXNwbGF5IHRoaXMgaGVscCB0ZXh0XG4iCiJcdC1hIC0t
YXNjaWlcdGRpc3BsYXkgdGhlIGRlY2ltYWwvb2N0YWwvaGV4IHZhbHVlcyBvZiB0aGUga2V5c1xu
IgoiXHQtcyAtLXNjYW5jb2Rlc1x0ZGlzcGxheSBvbmx5IHRoZSByYXcgc2Nhbi1jb2Rlc1xuIgoi
XHQtayAtLWtleWNvZGVzXHRkaXNwbGF5IG9ubHkgdGhlIGludGVycHJldGVkIGtleWNvZGVzIChk
ZWZhdWx0KVxuIgptc2dzdHIgIiIKInNob3drZXkgdmVyc2lvbiAlc1xuIgoiXG4iCiJhbnbkbmRu
aW5nOiBzaG93a2V5IFtmbGFnZ29yLi4uXVxuIgoiXG4iCiJ0aWxs5XRuYSBmbGFnZ29yIORyOlxu
IgoiXG4iCiJcdC1oIC0taGVscFx0dmlzYSBkZW4gaORyIGhq5GxwdGV4dGVuXG4iCiJcdC1hIC0t
YXNjaWlcdHZpc2EgZGVjaW1hbGEvb2t0YWxhL2hleGFkZWNpbWFsYSB25HJkZW4gZvZyIHRlY2tu
ZW5cbiIKIlx0LXMgLS1zY2FuY29kZXNcdHZpc2EgYmFyYSBkZSBy5WEgYXZs5HNuaW5nc2tvZGVy
bmFcbiIKIlx0LWsgLS1rZXljb2Rlc1x0dmlzYSBiYXJhIGRlIHRvbGthZGUgdGFuZ2VudGtvZGVy
bmEgKHN0YW5kYXJkdmFsKVxuIgoKIzogc3JjL3Nob3drZXkuYzoxNTcKbXNnaWQgIlxuUHJlc3Mg
YW55IGtleXMgLSBDdHJsLUQgd2lsbCB0ZXJtaW5hdGUgdGhpcyBwcm9ncmFtXG5cbiIKbXNnc3Ry
ICJcblRyeWNrIG7lZ29uIHRhbmdlbnQgLSBDdHJsLUQga29tbWVyIGF0dCBhdnNsdXRhIHByb2dy
YW1tZXRcblxuIgoKIzogc3JjL3Nob3drZXkuYzoyMjYKbXNnaWQgInByZXNzIGFueSBrZXkgKHBy
b2dyYW0gdGVybWluYXRlcyAxMHMgYWZ0ZXIgbGFzdCBrZXlwcmVzcykuLi5cbiIKbXNnc3RyICJ0
cnljayBu5WdvbiB0YW5nZW50IChwcm9ncmFtbWV0IGF2c2x1dGFzIDEwIHMgZWZ0ZXIgc2lzdGEg
dGFuZ2VudHRyeWNrbmluZykuLi5cbiIKCiM6IHNyYy9zaG93a2V5LmM6MjM0CiMsIGMtZm9ybWF0
Cm1zZ2lkICJrZXljb2RlICUzZCAlc1xuIgptc2dzdHIgInRhbmdlbnRrb2QgJTNkICVzXG4iCgoj
OiBzcmMvc2hvd2tleS5jOjIzNgptc2dpZCAicmVsZWFzZSIKbXNnc3RyICJzbORwcCIKCiM6IHNy
Yy9zaG93a2V5LmM6MjM3Cm1zZ2lkICJwcmVzcyIKbXNnc3RyICJ0cnljayIKCiM6IHNyYy92ZXJz
aW9uLmg6MTcKIywgYy1mb3JtYXQKbXNnaWQgIiVzIGZyb20gJXNcbiIKbXNnc3RyICIlcyBmcuVu
ICVzXG4iCg==
--=-=-=

                                The Translation Project robot, in the
                                name of your kind translation coordinator.
                                mailto:translation@iro.umontreal.ca

--=-=-=--

